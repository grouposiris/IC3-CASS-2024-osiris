magic
tech sky130A
magscale 1 2
timestamp 1731062359
<< obsli1 >>
rect 2760 2703 34316 34289
<< obsm1 >>
rect 14 2672 36786 34320
<< metal2 >>
rect 662 35678 718 36478
rect 1950 35678 2006 36478
rect 3238 35678 3294 36478
rect 4526 35678 4582 36478
rect 5814 35678 5870 36478
rect 7746 35678 7802 36478
rect 9034 35678 9090 36478
rect 10322 35678 10378 36478
rect 11610 35678 11666 36478
rect 12898 35678 12954 36478
rect 14186 35678 14242 36478
rect 15474 35678 15530 36478
rect 17406 35678 17462 36478
rect 18694 35678 18750 36478
rect 19982 35678 20038 36478
rect 21270 35678 21326 36478
rect 22558 35678 22614 36478
rect 23846 35678 23902 36478
rect 25134 35678 25190 36478
rect 26422 35678 26478 36478
rect 28354 35678 28410 36478
rect 29642 35678 29698 36478
rect 30930 35678 30986 36478
rect 32218 35678 32274 36478
rect 33506 35678 33562 36478
rect 34794 35678 34850 36478
rect 36082 35678 36138 36478
rect 18 0 74 800
rect 1306 0 1362 800
rect 2594 0 2650 800
rect 3882 0 3938 800
rect 5170 0 5226 800
rect 6458 0 6514 800
rect 7746 0 7802 800
rect 9034 0 9090 800
rect 10966 0 11022 800
rect 12254 0 12310 800
rect 13542 0 13598 800
rect 14830 0 14886 800
rect 16118 0 16174 800
rect 17406 0 17462 800
rect 18694 0 18750 800
rect 20626 0 20682 800
rect 21914 0 21970 800
rect 23202 0 23258 800
rect 24490 0 24546 800
rect 25778 0 25834 800
rect 27066 0 27122 800
rect 28354 0 28410 800
rect 29642 0 29698 800
rect 31574 0 31630 800
rect 32862 0 32918 800
rect 34150 0 34206 800
rect 35438 0 35494 800
rect 36726 0 36782 800
<< obsm2 >>
rect 20 35622 606 36145
rect 774 35622 1894 36145
rect 2062 35622 3182 36145
rect 3350 35622 4470 36145
rect 4638 35622 5758 36145
rect 5926 35622 7690 36145
rect 7858 35622 8978 36145
rect 9146 35622 10266 36145
rect 10434 35622 11554 36145
rect 11722 35622 12842 36145
rect 13010 35622 14130 36145
rect 14298 35622 15418 36145
rect 15586 35622 17350 36145
rect 17518 35622 18638 36145
rect 18806 35622 19926 36145
rect 20094 35622 21214 36145
rect 21382 35622 22502 36145
rect 22670 35622 23790 36145
rect 23958 35622 25078 36145
rect 25246 35622 26366 36145
rect 26534 35622 28298 36145
rect 28466 35622 29586 36145
rect 29754 35622 30874 36145
rect 31042 35622 32162 36145
rect 32330 35622 33450 36145
rect 33618 35622 34738 36145
rect 34906 35622 36026 36145
rect 36194 35622 36780 36145
rect 20 856 36780 35622
rect 130 800 1250 856
rect 1418 800 2538 856
rect 2706 800 3826 856
rect 3994 800 5114 856
rect 5282 800 6402 856
rect 6570 800 7690 856
rect 7858 800 8978 856
rect 9146 800 10910 856
rect 11078 800 12198 856
rect 12366 800 13486 856
rect 13654 800 14774 856
rect 14942 800 16062 856
rect 16230 800 17350 856
rect 17518 800 18638 856
rect 18806 800 20570 856
rect 20738 800 21858 856
rect 22026 800 23146 856
rect 23314 800 24434 856
rect 24602 800 25722 856
rect 25890 800 27010 856
rect 27178 800 28298 856
rect 28466 800 29586 856
rect 29754 800 31518 856
rect 31686 800 32806 856
rect 32974 800 34094 856
rect 34262 800 35382 856
rect 35550 800 36670 856
<< metal3 >>
rect 0 36048 800 36168
rect 36302 35368 37102 35488
rect 0 34688 800 34808
rect 36302 34008 37102 34128
rect 0 33328 800 33448
rect 36302 32648 37102 32768
rect 0 31288 800 31408
rect 36302 31288 37102 31408
rect 0 29928 800 30048
rect 36302 29928 37102 30048
rect 0 28568 800 28688
rect 36302 28568 37102 28688
rect 0 27208 800 27328
rect 36302 27208 37102 27328
rect 0 25848 800 25968
rect 36302 25848 37102 25968
rect 0 24488 800 24608
rect 36302 23808 37102 23928
rect 0 23128 800 23248
rect 36302 22448 37102 22568
rect 0 21088 800 21208
rect 36302 21088 37102 21208
rect 0 19728 800 19848
rect 36302 19728 37102 19848
rect 0 18368 800 18488
rect 36302 18368 37102 18488
rect 0 17008 800 17128
rect 36302 17008 37102 17128
rect 0 15648 800 15768
rect 36302 15648 37102 15768
rect 0 14288 800 14408
rect 36302 13608 37102 13728
rect 0 12928 800 13048
rect 36302 12248 37102 12368
rect 0 11568 800 11688
rect 36302 10888 37102 11008
rect 0 9528 800 9648
rect 36302 9528 37102 9648
rect 0 8168 800 8288
rect 36302 8168 37102 8288
rect 0 6808 800 6928
rect 36302 6808 37102 6928
rect 0 5448 800 5568
rect 36302 5448 37102 5568
rect 0 4088 800 4208
rect 36302 4088 37102 4208
rect 0 2728 800 2848
rect 36302 2048 37102 2168
rect 0 1368 800 1488
rect 36302 688 37102 808
<< obsm3 >>
rect 880 35968 36302 36141
rect 800 35568 36302 35968
rect 800 35288 36222 35568
rect 800 34888 36302 35288
rect 880 34608 36302 34888
rect 800 34208 36302 34608
rect 800 33928 36222 34208
rect 800 33528 36302 33928
rect 880 33248 36302 33528
rect 800 32848 36302 33248
rect 800 32568 36222 32848
rect 800 31488 36302 32568
rect 880 31208 36222 31488
rect 800 30128 36302 31208
rect 880 29848 36222 30128
rect 800 28768 36302 29848
rect 880 28488 36222 28768
rect 800 27408 36302 28488
rect 880 27128 36222 27408
rect 800 26048 36302 27128
rect 880 25768 36222 26048
rect 800 24688 36302 25768
rect 880 24408 36302 24688
rect 800 24008 36302 24408
rect 800 23728 36222 24008
rect 800 23328 36302 23728
rect 880 23048 36302 23328
rect 800 22648 36302 23048
rect 800 22368 36222 22648
rect 800 21288 36302 22368
rect 880 21008 36222 21288
rect 800 19928 36302 21008
rect 880 19648 36222 19928
rect 800 18568 36302 19648
rect 880 18288 36222 18568
rect 800 17208 36302 18288
rect 880 16928 36222 17208
rect 800 15848 36302 16928
rect 880 15568 36222 15848
rect 800 14488 36302 15568
rect 880 14208 36302 14488
rect 800 13808 36302 14208
rect 800 13528 36222 13808
rect 800 13128 36302 13528
rect 880 12848 36302 13128
rect 800 12448 36302 12848
rect 800 12168 36222 12448
rect 800 11768 36302 12168
rect 880 11488 36302 11768
rect 800 11088 36302 11488
rect 800 10808 36222 11088
rect 800 9728 36302 10808
rect 880 9448 36222 9728
rect 800 8368 36302 9448
rect 880 8088 36222 8368
rect 800 7008 36302 8088
rect 880 6728 36222 7008
rect 800 5648 36302 6728
rect 880 5368 36222 5648
rect 800 4288 36302 5368
rect 880 4008 36222 4288
rect 800 2928 36302 4008
rect 880 2648 36302 2928
rect 800 2248 36302 2648
rect 800 1968 36222 2248
rect 800 1568 36302 1968
rect 880 1288 36302 1568
rect 800 888 36302 1288
rect 800 718 36222 888
<< metal4 >>
rect 6544 2672 6864 34320
rect 7204 2672 7524 34320
rect 14433 2672 14753 34320
rect 15093 2672 15413 34320
rect 22322 2672 22642 34320
rect 22982 2672 23302 34320
rect 30211 2672 30531 34320
rect 30871 2672 31191 34320
<< obsm4 >>
rect 5579 3027 6464 33285
rect 6944 3027 7124 33285
rect 7604 3027 14353 33285
rect 14833 3027 15013 33285
rect 15493 3027 22242 33285
rect 22722 3027 22902 33285
rect 23382 3027 27909 33285
<< labels >>
rlabel metal2 s 11610 35678 11666 36478 6 clk
port 1 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 i_start_rx
port 2 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 i_uart_rx
port 3 nsew signal input
rlabel metal2 s 19982 35678 20038 36478 6 o_uart_tx
port 4 nsew signal output
rlabel metal3 s 0 34688 800 34808 6 rst
port 5 nsew signal input
rlabel metal4 s 6544 2672 6864 34320 6 vccd1
port 6 nsew power bidirectional
rlabel metal4 s 14433 2672 14753 34320 6 vccd1
port 6 nsew power bidirectional
rlabel metal4 s 22322 2672 22642 34320 6 vccd1
port 6 nsew power bidirectional
rlabel metal4 s 30211 2672 30531 34320 6 vccd1
port 6 nsew power bidirectional
rlabel metal4 s 7204 2672 7524 34320 6 vssd1
port 7 nsew ground bidirectional
rlabel metal4 s 15093 2672 15413 34320 6 vssd1
port 7 nsew ground bidirectional
rlabel metal4 s 22982 2672 23302 34320 6 vssd1
port 7 nsew ground bidirectional
rlabel metal4 s 30871 2672 31191 34320 6 vssd1
port 7 nsew ground bidirectional
rlabel metal3 s 36302 12248 37102 12368 6 wb_ack_i
port 8 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 wb_adr_o[0]
port 9 nsew signal output
rlabel metal2 s 23846 35678 23902 36478 6 wb_adr_o[10]
port 10 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 wb_adr_o[11]
port 11 nsew signal output
rlabel metal3 s 0 12928 800 13048 6 wb_adr_o[12]
port 12 nsew signal output
rlabel metal3 s 36302 28568 37102 28688 6 wb_adr_o[13]
port 13 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 wb_adr_o[14]
port 14 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 wb_adr_o[15]
port 15 nsew signal output
rlabel metal3 s 36302 6808 37102 6928 6 wb_adr_o[16]
port 16 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 wb_adr_o[17]
port 17 nsew signal output
rlabel metal3 s 36302 18368 37102 18488 6 wb_adr_o[18]
port 18 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 wb_adr_o[19]
port 19 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 wb_adr_o[1]
port 20 nsew signal output
rlabel metal2 s 32218 35678 32274 36478 6 wb_adr_o[20]
port 21 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 wb_adr_o[21]
port 22 nsew signal output
rlabel metal3 s 36302 5448 37102 5568 6 wb_adr_o[22]
port 23 nsew signal output
rlabel metal3 s 36302 19728 37102 19848 6 wb_adr_o[23]
port 24 nsew signal output
rlabel metal3 s 36302 32648 37102 32768 6 wb_adr_o[24]
port 25 nsew signal output
rlabel metal2 s 4526 35678 4582 36478 6 wb_adr_o[25]
port 26 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 wb_adr_o[26]
port 27 nsew signal output
rlabel metal2 s 26422 35678 26478 36478 6 wb_adr_o[27]
port 28 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 wb_adr_o[28]
port 29 nsew signal output
rlabel metal2 s 34794 35678 34850 36478 6 wb_adr_o[29]
port 30 nsew signal output
rlabel metal3 s 36302 34008 37102 34128 6 wb_adr_o[2]
port 31 nsew signal output
rlabel metal2 s 7746 0 7802 800 6 wb_adr_o[30]
port 32 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 wb_adr_o[31]
port 33 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 wb_adr_o[3]
port 34 nsew signal output
rlabel metal3 s 36302 35368 37102 35488 6 wb_adr_o[4]
port 35 nsew signal output
rlabel metal2 s 30930 35678 30986 36478 6 wb_adr_o[5]
port 36 nsew signal output
rlabel metal3 s 36302 688 37102 808 6 wb_adr_o[6]
port 37 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 wb_adr_o[7]
port 38 nsew signal output
rlabel metal3 s 36302 15648 37102 15768 6 wb_adr_o[8]
port 39 nsew signal output
rlabel metal3 s 36302 10888 37102 11008 6 wb_adr_o[9]
port 40 nsew signal output
rlabel metal2 s 12898 35678 12954 36478 6 wb_cyc_o
port 41 nsew signal output
rlabel metal2 s 14186 35678 14242 36478 6 wb_dat_i[0]
port 42 nsew signal input
rlabel metal3 s 36302 27208 37102 27328 6 wb_dat_i[10]
port 43 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 wb_dat_i[11]
port 44 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 wb_dat_i[12]
port 45 nsew signal input
rlabel metal3 s 36302 29928 37102 30048 6 wb_dat_i[13]
port 46 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 wb_dat_i[14]
port 47 nsew signal input
rlabel metal2 s 21270 35678 21326 36478 6 wb_dat_i[15]
port 48 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 wb_dat_i[16]
port 49 nsew signal input
rlabel metal2 s 10322 35678 10378 36478 6 wb_dat_i[17]
port 50 nsew signal input
rlabel metal2 s 15474 35678 15530 36478 6 wb_dat_i[18]
port 51 nsew signal input
rlabel metal3 s 36302 31288 37102 31408 6 wb_dat_i[19]
port 52 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 wb_dat_i[1]
port 53 nsew signal input
rlabel metal2 s 18694 35678 18750 36478 6 wb_dat_i[20]
port 54 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 wb_dat_i[21]
port 55 nsew signal input
rlabel metal3 s 36302 8168 37102 8288 6 wb_dat_i[22]
port 56 nsew signal input
rlabel metal3 s 36302 22448 37102 22568 6 wb_dat_i[23]
port 57 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 wb_dat_i[24]
port 58 nsew signal input
rlabel metal2 s 22558 35678 22614 36478 6 wb_dat_i[25]
port 59 nsew signal input
rlabel metal2 s 7746 35678 7802 36478 6 wb_dat_i[26]
port 60 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 wb_dat_i[27]
port 61 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 wb_dat_i[28]
port 62 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 wb_dat_i[29]
port 63 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wb_dat_i[2]
port 64 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 wb_dat_i[30]
port 65 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 wb_dat_i[31]
port 66 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 wb_dat_i[3]
port 67 nsew signal input
rlabel metal3 s 36302 9528 37102 9648 6 wb_dat_i[4]
port 68 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 wb_dat_i[5]
port 69 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 wb_dat_i[6]
port 70 nsew signal input
rlabel metal3 s 36302 2048 37102 2168 6 wb_dat_i[7]
port 71 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 wb_dat_i[8]
port 72 nsew signal input
rlabel metal3 s 36302 13608 37102 13728 6 wb_dat_i[9]
port 73 nsew signal input
rlabel metal3 s 36302 23808 37102 23928 6 wb_dat_o[0]
port 74 nsew signal output
rlabel metal2 s 29642 0 29698 800 6 wb_dat_o[10]
port 75 nsew signal output
rlabel metal3 s 36302 25848 37102 25968 6 wb_dat_o[11]
port 76 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 wb_dat_o[12]
port 77 nsew signal output
rlabel metal2 s 662 35678 718 36478 6 wb_dat_o[13]
port 78 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 wb_dat_o[14]
port 79 nsew signal output
rlabel metal2 s 18 0 74 800 6 wb_dat_o[15]
port 80 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 wb_dat_o[16]
port 81 nsew signal output
rlabel metal2 s 5814 35678 5870 36478 6 wb_dat_o[17]
port 82 nsew signal output
rlabel metal2 s 17406 35678 17462 36478 6 wb_dat_o[18]
port 83 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 wb_dat_o[19]
port 84 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 wb_dat_o[1]
port 85 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 wb_dat_o[20]
port 86 nsew signal output
rlabel metal2 s 1306 0 1362 800 6 wb_dat_o[21]
port 87 nsew signal output
rlabel metal2 s 33506 35678 33562 36478 6 wb_dat_o[22]
port 88 nsew signal output
rlabel metal2 s 25134 35678 25190 36478 6 wb_dat_o[23]
port 89 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 wb_dat_o[24]
port 90 nsew signal output
rlabel metal2 s 36082 35678 36138 36478 6 wb_dat_o[25]
port 91 nsew signal output
rlabel metal3 s 36302 4088 37102 4208 6 wb_dat_o[26]
port 92 nsew signal output
rlabel metal2 s 1950 35678 2006 36478 6 wb_dat_o[27]
port 93 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 wb_dat_o[28]
port 94 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 wb_dat_o[29]
port 95 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 wb_dat_o[2]
port 96 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 wb_dat_o[30]
port 97 nsew signal output
rlabel metal3 s 36302 21088 37102 21208 6 wb_dat_o[31]
port 98 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 wb_dat_o[3]
port 99 nsew signal output
rlabel metal2 s 29642 35678 29698 36478 6 wb_dat_o[4]
port 100 nsew signal output
rlabel metal2 s 28354 35678 28410 36478 6 wb_dat_o[5]
port 101 nsew signal output
rlabel metal2 s 3238 35678 3294 36478 6 wb_dat_o[6]
port 102 nsew signal output
rlabel metal2 s 9034 35678 9090 36478 6 wb_dat_o[7]
port 103 nsew signal output
rlabel metal2 s 24490 0 24546 800 6 wb_dat_o[8]
port 104 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 wb_dat_o[9]
port 105 nsew signal output
rlabel metal3 s 0 33328 800 33448 6 wb_stb_o
port 106 nsew signal output
rlabel metal3 s 36302 17008 37102 17128 6 wb_we_o
port 107 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 37102 36478
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3955736
string GDS_FILE /home/roliveira/Desktop/osiris_i/openlane/uart_wbs_bridge/runs/oeb_fix/results/signoff/uart_wbs_bridge.magic.gds
string GDS_START 561540
<< end >>

