magic
tech sky130A
magscale 1 2
timestamp 1731186435
<< obsli1 >>
rect 7360 2703 282164 308465
<< obsm1 >>
rect 14 2672 282886 308496
<< metal2 >>
rect 6458 310200 6514 311000
rect 49606 310200 49662 311000
rect 92754 310200 92810 311000
rect 135902 310200 135958 311000
rect 179050 310200 179106 311000
rect 222198 310200 222254 311000
rect 265346 310200 265402 311000
rect 18 0 74 800
rect 42522 0 42578 800
rect 85670 0 85726 800
rect 128818 0 128874 800
rect 171966 0 172022 800
rect 215114 0 215170 800
rect 258262 0 258318 800
<< obsm2 >>
rect 20 310144 6402 310298
rect 6570 310144 49550 310298
rect 49718 310144 92698 310298
rect 92866 310144 135846 310298
rect 136014 310144 178994 310298
rect 179162 310144 222142 310298
rect 222310 310144 265290 310298
rect 265458 310144 282882 310298
rect 20 856 282882 310144
rect 130 800 42466 856
rect 42634 800 85614 856
rect 85782 800 128762 856
rect 128930 800 171910 856
rect 172078 800 215058 856
rect 215226 800 258206 856
rect 258374 800 282882 856
<< metal3 >>
rect 286000 288328 286800 288448
rect 0 272688 800 272808
rect 286000 242768 286800 242888
rect 0 227128 800 227248
rect 286000 197208 286800 197328
rect 0 181568 800 181688
rect 286000 151648 286800 151768
rect 0 136008 800 136128
rect 286000 106088 286800 106208
rect 0 90448 800 90568
rect 286000 60528 286800 60648
rect 0 44888 800 45008
rect 286000 14968 286800 15088
<< obsm3 >>
rect 800 288528 286000 308481
rect 800 288248 285920 288528
rect 800 272888 286000 288248
rect 880 272608 286000 272888
rect 800 242968 286000 272608
rect 800 242688 285920 242968
rect 800 227328 286000 242688
rect 880 227048 286000 227328
rect 800 197408 286000 227048
rect 800 197128 285920 197408
rect 800 181768 286000 197128
rect 880 181488 286000 181768
rect 800 151848 286000 181488
rect 800 151568 285920 151848
rect 800 136208 286000 151568
rect 880 135928 286000 136208
rect 800 106288 286000 135928
rect 800 106008 285920 106288
rect 800 90648 286000 106008
rect 880 90368 286000 90648
rect 800 60728 286000 90368
rect 800 60448 285920 60728
rect 800 45088 286000 60448
rect 880 44808 286000 45088
rect 800 15168 286000 44808
rect 800 14888 285920 15168
rect 800 2687 286000 14888
<< metal4 >>
rect 5180 540 5500 310628
rect 5840 1200 6160 309968
rect 10464 540 10784 310628
rect 11124 540 11444 310628
rect 41184 294877 41504 310628
rect 41844 294877 42164 310628
rect 71904 294877 72224 310628
rect 72564 294877 72884 310628
rect 102624 294877 102944 310628
rect 103284 294877 103604 310628
rect 133344 294877 133664 310628
rect 134004 294877 134324 310628
rect 164064 294877 164384 310628
rect 164724 294877 165044 310628
rect 41184 144677 41504 161371
rect 41844 144677 42164 161371
rect 71904 144677 72224 161371
rect 72564 144677 72884 161371
rect 102624 144677 102944 161371
rect 103284 144677 103604 161371
rect 133344 144677 133664 161371
rect 134004 144677 134324 161371
rect 164064 144677 164384 161371
rect 164724 144677 165044 161371
rect 179516 160432 179836 238864
rect 180252 160432 180572 238864
rect 179516 103312 179836 145840
rect 180252 103312 180572 145840
rect 41184 540 41504 11171
rect 41844 540 42164 11171
rect 71904 540 72224 11171
rect 72564 540 72884 11171
rect 102624 540 102944 11171
rect 103284 540 103604 11171
rect 133344 540 133664 11171
rect 134004 540 134324 11171
rect 164064 540 164384 11171
rect 164724 540 165044 11171
rect 194784 540 195104 310628
rect 195444 540 195764 310628
rect 225504 235093 225824 310628
rect 226164 235093 226484 310628
rect 225504 69911 225824 106619
rect 226164 69911 226484 106619
rect 225504 540 225824 35413
rect 226164 540 226484 35413
rect 256224 540 256544 310628
rect 256884 540 257204 310628
rect 276668 103312 276988 238864
rect 277404 103312 277724 238864
rect 283364 1200 283684 309968
rect 284024 540 284344 310628
<< obsm4 >>
rect 21472 238944 194704 293181
rect 21472 161451 179436 238944
rect 21472 144597 41104 161451
rect 41584 144597 41764 161451
rect 42244 144597 71824 161451
rect 72304 144597 72484 161451
rect 72964 144597 102544 161451
rect 103024 144597 103204 161451
rect 103684 144597 133264 161451
rect 133744 144597 133924 161451
rect 134404 144597 163984 161451
rect 164464 144597 164644 161451
rect 165124 160352 179436 161451
rect 179916 160352 180172 238944
rect 180652 160352 194704 238944
rect 165124 145920 194704 160352
rect 165124 144597 179436 145920
rect 21472 103232 179436 144597
rect 179916 103232 180172 145920
rect 180652 103232 194704 145920
rect 21472 12275 194704 103232
rect 195184 12275 195364 293181
rect 195844 235013 225424 293181
rect 225904 235013 226084 293181
rect 226564 235013 256144 293181
rect 195844 106699 256144 235013
rect 195844 69831 225424 106699
rect 225904 69831 226084 106699
rect 226564 69831 256144 106699
rect 195844 35493 256144 69831
rect 195844 12275 225424 35493
rect 225904 12275 226084 35493
rect 226564 12275 256144 35493
rect 256624 12275 256804 293181
rect 257284 12275 272629 293181
<< metal5 >>
rect 5180 310308 284344 310628
rect 5840 309648 283684 309968
rect 5180 282274 284344 282594
rect 5180 281614 284344 281934
rect 5180 251638 284344 251958
rect 5180 250978 284344 251298
rect 5180 221002 284344 221322
rect 5180 220342 284344 220662
rect 5180 190366 284344 190686
rect 5180 189706 284344 190026
rect 5180 159730 284344 160050
rect 5180 159070 284344 159390
rect 5180 129094 284344 129414
rect 5180 128434 284344 128754
rect 5180 98458 284344 98778
rect 5180 97798 284344 98118
rect 5180 67822 284344 68142
rect 5180 67162 284344 67482
rect 5180 37186 284344 37506
rect 5180 36526 284344 36846
rect 5180 6550 284344 6870
rect 5180 5890 284344 6210
rect 5840 1200 283684 1520
rect 5180 540 284344 860
<< labels >>
rlabel metal3 s 286000 14968 286800 15088 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 286000 106088 286800 106208 6 io_in[1]
port 2 nsew signal input
rlabel metal2 s 128818 0 128874 800 6 io_in[2]
port 3 nsew signal input
rlabel metal3 s 0 227128 800 227248 6 io_in[3]
port 4 nsew signal input
rlabel metal3 s 0 90448 800 90568 6 io_in[4]
port 5 nsew signal input
rlabel metal3 s 0 272688 800 272808 6 io_oeb[0]
port 6 nsew signal output
rlabel metal2 s 265346 310200 265402 311000 6 io_oeb[10]
port 7 nsew signal output
rlabel metal2 s 215114 0 215170 800 6 io_oeb[11]
port 8 nsew signal output
rlabel metal3 s 0 44888 800 45008 6 io_oeb[1]
port 9 nsew signal output
rlabel metal2 s 222198 310200 222254 311000 6 io_oeb[2]
port 10 nsew signal output
rlabel metal3 s 286000 288328 286800 288448 6 io_oeb[3]
port 11 nsew signal output
rlabel metal3 s 0 136008 800 136128 6 io_oeb[4]
port 12 nsew signal output
rlabel metal2 s 49606 310200 49662 311000 6 io_oeb[5]
port 13 nsew signal output
rlabel metal2 s 258262 0 258318 800 6 io_oeb[6]
port 14 nsew signal output
rlabel metal2 s 18 0 74 800 6 io_oeb[7]
port 15 nsew signal output
rlabel metal2 s 42522 0 42578 800 6 io_oeb[8]
port 16 nsew signal output
rlabel metal2 s 92754 310200 92810 311000 6 io_oeb[9]
port 17 nsew signal output
rlabel metal3 s 286000 60528 286800 60648 6 io_out[0]
port 18 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 io_out[1]
port 19 nsew signal output
rlabel metal3 s 286000 197208 286800 197328 6 io_out[2]
port 20 nsew signal output
rlabel metal3 s 286000 242768 286800 242888 6 io_out[3]
port 21 nsew signal output
rlabel metal2 s 135902 310200 135958 311000 6 io_out[4]
port 22 nsew signal output
rlabel metal2 s 179050 310200 179106 311000 6 io_out[5]
port 23 nsew signal output
rlabel metal2 s 171966 0 172022 800 6 io_out[6]
port 24 nsew signal output
rlabel metal3 s 0 181568 800 181688 6 io_out[7]
port 25 nsew signal output
rlabel metal2 s 6458 310200 6514 311000 6 io_out[8]
port 26 nsew signal output
rlabel metal4 s 5840 1200 6160 309968 6 vccd1
port 27 nsew power bidirectional
rlabel metal5 s 5840 1200 283684 1520 6 vccd1
port 27 nsew power bidirectional
rlabel metal5 s 5840 309648 283684 309968 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 283364 1200 283684 309968 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 10464 540 10784 310628 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 41184 540 41504 11171 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 41184 144677 41504 161371 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 41184 294877 41504 310628 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 71904 540 72224 11171 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 71904 144677 72224 161371 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 71904 294877 72224 310628 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 102624 540 102944 11171 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 102624 144677 102944 161371 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 102624 294877 102944 310628 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 133344 540 133664 11171 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 133344 144677 133664 161371 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 133344 294877 133664 310628 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 164064 540 164384 11171 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 164064 144677 164384 161371 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 164064 294877 164384 310628 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 194784 540 195104 310628 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 225504 540 225824 35413 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 225504 69911 225824 106619 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 225504 235093 225824 310628 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 256224 540 256544 310628 6 vccd1
port 27 nsew power bidirectional
rlabel metal5 s 5180 5890 284344 6210 6 vccd1
port 27 nsew power bidirectional
rlabel metal5 s 5180 36526 284344 36846 6 vccd1
port 27 nsew power bidirectional
rlabel metal5 s 5180 67162 284344 67482 6 vccd1
port 27 nsew power bidirectional
rlabel metal5 s 5180 97798 284344 98118 6 vccd1
port 27 nsew power bidirectional
rlabel metal5 s 5180 128434 284344 128754 6 vccd1
port 27 nsew power bidirectional
rlabel metal5 s 5180 159070 284344 159390 6 vccd1
port 27 nsew power bidirectional
rlabel metal5 s 5180 189706 284344 190026 6 vccd1
port 27 nsew power bidirectional
rlabel metal5 s 5180 220342 284344 220662 6 vccd1
port 27 nsew power bidirectional
rlabel metal5 s 5180 250978 284344 251298 6 vccd1
port 27 nsew power bidirectional
rlabel metal5 s 5180 281614 284344 281934 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 179516 103312 179836 145840 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 179516 160432 179836 238864 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 276668 103312 276988 238864 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 5180 540 5500 310628 6 vssd1
port 28 nsew ground bidirectional
rlabel metal5 s 5180 540 284344 860 6 vssd1
port 28 nsew ground bidirectional
rlabel metal5 s 5180 310308 284344 310628 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 284024 540 284344 310628 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 11124 540 11444 310628 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 41844 540 42164 11171 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 41844 144677 42164 161371 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 41844 294877 42164 310628 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 72564 540 72884 11171 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 72564 144677 72884 161371 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 72564 294877 72884 310628 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 103284 540 103604 11171 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 103284 144677 103604 161371 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 103284 294877 103604 310628 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 134004 540 134324 11171 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 134004 144677 134324 161371 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 134004 294877 134324 310628 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 164724 540 165044 11171 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 164724 144677 165044 161371 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 164724 294877 165044 310628 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 195444 540 195764 310628 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 226164 540 226484 35413 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 226164 69911 226484 106619 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 226164 235093 226484 310628 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 256884 540 257204 310628 6 vssd1
port 28 nsew ground bidirectional
rlabel metal5 s 5180 6550 284344 6870 6 vssd1
port 28 nsew ground bidirectional
rlabel metal5 s 5180 37186 284344 37506 6 vssd1
port 28 nsew ground bidirectional
rlabel metal5 s 5180 67822 284344 68142 6 vssd1
port 28 nsew ground bidirectional
rlabel metal5 s 5180 98458 284344 98778 6 vssd1
port 28 nsew ground bidirectional
rlabel metal5 s 5180 129094 284344 129414 6 vssd1
port 28 nsew ground bidirectional
rlabel metal5 s 5180 159730 284344 160050 6 vssd1
port 28 nsew ground bidirectional
rlabel metal5 s 5180 190366 284344 190686 6 vssd1
port 28 nsew ground bidirectional
rlabel metal5 s 5180 221002 284344 221322 6 vssd1
port 28 nsew ground bidirectional
rlabel metal5 s 5180 251638 284344 251958 6 vssd1
port 28 nsew ground bidirectional
rlabel metal5 s 5180 282274 284344 282594 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 180252 103312 180572 145840 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 180252 160432 180572 238864 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 277404 103312 277724 238864 6 vssd1
port 28 nsew ground bidirectional
rlabel metal3 s 286000 151648 286800 151768 6 wb_clk_i
port 29 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 286800 311000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 131596944
string GDS_FILE /home/roliveira/Desktop/osiris_i/openlane/osiris_i_wrapper/runs/lvs/results/signoff/osiris_i_wrapper.magic.gds
string GDS_START 110134570
<< end >>

