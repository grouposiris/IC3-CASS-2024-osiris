* NGSPICE file created from uart_wbs_bridge.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

.subckt uart_wbs_bridge clk i_start_rx i_uart_rx o_uart_tx rst vccd1 vssd1 wb_ack_i
+ wb_adr_o[0] wb_adr_o[10] wb_adr_o[11] wb_adr_o[12] wb_adr_o[13] wb_adr_o[14] wb_adr_o[15]
+ wb_adr_o[16] wb_adr_o[17] wb_adr_o[18] wb_adr_o[19] wb_adr_o[1] wb_adr_o[20] wb_adr_o[21]
+ wb_adr_o[22] wb_adr_o[23] wb_adr_o[24] wb_adr_o[25] wb_adr_o[26] wb_adr_o[27] wb_adr_o[28]
+ wb_adr_o[29] wb_adr_o[2] wb_adr_o[30] wb_adr_o[31] wb_adr_o[3] wb_adr_o[4] wb_adr_o[5]
+ wb_adr_o[6] wb_adr_o[7] wb_adr_o[8] wb_adr_o[9] wb_cyc_o wb_dat_i[0] wb_dat_i[10]
+ wb_dat_i[11] wb_dat_i[12] wb_dat_i[13] wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17]
+ wb_dat_i[18] wb_dat_i[19] wb_dat_i[1] wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23]
+ wb_dat_i[24] wb_dat_i[25] wb_dat_i[26] wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2]
+ wb_dat_i[30] wb_dat_i[31] wb_dat_i[3] wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7]
+ wb_dat_i[8] wb_dat_i[9] wb_dat_o[0] wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13]
+ wb_dat_o[14] wb_dat_o[15] wb_dat_o[16] wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1]
+ wb_dat_o[20] wb_dat_o[21] wb_dat_o[22] wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26]
+ wb_dat_o[27] wb_dat_o[28] wb_dat_o[29] wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3]
+ wb_dat_o[4] wb_dat_o[5] wb_dat_o[6] wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_stb_o
+ wb_we_o
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold351 _0845_/X vssd1 vssd1 vccd1 vccd1 _1608_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold362 _1613_/Q vssd1 vssd1 vccd1 vccd1 _0798_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold340 _1615_/Q vssd1 vssd1 vccd1 vccd1 _0828_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold373 _1588_/Q vssd1 vssd1 vccd1 vccd1 hold373/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 _1585_/Q vssd1 vssd1 vccd1 vccd1 hold54/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1270_ _1402_/A vssd1 vssd1 vccd1 vccd1 _1270_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_46_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1606_ _1625_/CLK _1606_/D _1388_/Y vssd1 vssd1 vccd1 vccd1 _1606_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_1_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0985_ _1100_/A _1100_/C _1192_/C vssd1 vssd1 vccd1 vccd1 _1027_/A sky130_fd_sc_hd__or3b_1
X_1537_ _1548_/CLK _1537_/D _1319_/Y vssd1 vssd1 vccd1 vccd1 _1537_/Q sky130_fd_sc_hd__dfrtp_1
X_1399_ _1409_/A vssd1 vssd1 vccd1 vccd1 _1399_/Y sky130_fd_sc_hd__inv_2
Xfanout127 _1416_/A vssd1 vssd1 vccd1 vccd1 _1384_/A sky130_fd_sc_hd__buf_8
X_1468_ _1605_/CLK _1468_/D _1250_/Y vssd1 vssd1 vccd1 vccd1 _1468_/Q sky130_fd_sc_hd__dfrtp_1
Xfanout116 hold80/X vssd1 vssd1 vccd1 vccd1 _1100_/B sky130_fd_sc_hd__clkbuf_8
Xfanout105 _1173_/S vssd1 vssd1 vccd1 vccd1 _1168_/S sky130_fd_sc_hd__buf_6
XFILLER_0_49_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold181 _1457_/Q vssd1 vssd1 vccd1 vccd1 hold181/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 _0765_/X vssd1 vssd1 vccd1 vccd1 _1628_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold170 _1133_/X vssd1 vssd1 vccd1 vccd1 _1458_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0770_ _1623_/Q _1622_/Q _0795_/B _1608_/Q vssd1 vssd1 vccd1 vccd1 _0773_/B sky130_fd_sc_hd__or4bb_1
X_1322_ _1387_/A vssd1 vssd1 vccd1 vccd1 _1322_/Y sky130_fd_sc_hd__inv_2
X_1253_ _1339_/A vssd1 vssd1 vccd1 vccd1 _1253_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1106__A0 _0995_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1113__S _1135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1184_ _1184_/A _1184_/B vssd1 vssd1 vccd1 vccd1 _1185_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_54_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0968_ _1140_/A _1073_/B vssd1 vssd1 vccd1 vccd1 _1068_/S sky130_fd_sc_hd__nand2_2
XFILLER_0_19_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0899_ input1/X _0933_/B vssd1 vssd1 vccd1 vccd1 _0925_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_40_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0822_ _0822_/A _0836_/A vssd1 vssd1 vccd1 vccd1 _0822_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_24_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1108__S _1135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0753_ _0753_/A _1584_/Q _0764_/B _0753_/D vssd1 vssd1 vccd1 vccd1 _0753_/X sky130_fd_sc_hd__or4_1
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1305_ _1404_/A vssd1 vssd1 vccd1 vccd1 _1305_/Y sky130_fd_sc_hd__inv_2
X_1236_ _1339_/A vssd1 vssd1 vccd1 vccd1 _1236_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_19_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1098_ _1098_/A _1098_/B vssd1 vssd1 vccd1 vccd1 _1098_/X sky130_fd_sc_hd__and2_1
X_1167_ hold36/X _1430_/Q _1168_/S vssd1 vssd1 vccd1 vccd1 hold37/A sky130_fd_sc_hd__mux2_1
XFILLER_0_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1088__A2 input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1021_ _1021_/A _1027_/B vssd1 vssd1 vccd1 vccd1 _1021_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_56_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0805_ _0813_/A _0813_/B vssd1 vssd1 vccd1 vccd1 _0805_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_16_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0736_ _0917_/A _0741_/B _0741_/C _0736_/D vssd1 vssd1 vccd1 vccd1 _0753_/D sky130_fd_sc_hd__or4_4
XANTENNA__1012__A2 _1059_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1219_ _1397_/A vssd1 vssd1 vccd1 vccd1 _1219_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_47_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold52 hold52/A vssd1 vssd1 vccd1 vccd1 hold52/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold74 hold74/A vssd1 vssd1 vccd1 vccd1 hold74/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 hold63/A vssd1 vssd1 vccd1 vccd1 hold63/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_42_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold85 hold85/A vssd1 vssd1 vccd1 vccd1 hold85/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 hold96/A vssd1 vssd1 vccd1 vccd1 hold96/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1570_ _1583_/CLK _1570_/D _1352_/Y vssd1 vssd1 vccd1 vccd1 _1570_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1004_ _0981_/A _1100_/C _1192_/B vssd1 vssd1 vccd1 vccd1 _1005_/B sky130_fd_sc_hd__and3b_1
XANTENNA__1121__S _1133_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0719_ _0967_/B vssd1 vssd1 vccd1 vccd1 _1141_/B sky130_fd_sc_hd__inv_2
XFILLER_0_50_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput75 _1469_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[13] sky130_fd_sc_hd__buf_12
Xoutput64 _1428_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[4] sky130_fd_sc_hd__buf_12
XFILLER_0_50_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput42 _1437_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[13] sky130_fd_sc_hd__buf_12
Xoutput53 _1447_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[23] sky130_fd_sc_hd__buf_12
Xoutput97 _1460_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[4] sky130_fd_sc_hd__buf_12
Xoutput86 _1479_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[23] sky130_fd_sc_hd__buf_12
XFILLER_0_53_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0974__B2 _1059_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1622_ _1623_/CLK _1622_/D _1404_/Y vssd1 vssd1 vccd1 vccd1 _1622_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1484_ _1632_/CLK _1484_/D _1266_/Y vssd1 vssd1 vccd1 vccd1 _1484_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1553_ _1600_/CLK _1553_/D _1335_/Y vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__dfrtp_1
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1116__S _1133_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold385 _1529_/Q vssd1 vssd1 vccd1 vccd1 hold385/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 _0829_/X vssd1 vssd1 vccd1 vccd1 _0830_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold352 _1622_/Q vssd1 vssd1 vccd1 vccd1 _0807_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold374 _1594_/Q vssd1 vssd1 vccd1 vccd1 hold374/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold363 _1419_/Q vssd1 vssd1 vccd1 vccd1 hold363/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold330 _1418_/Q vssd1 vssd1 vccd1 vccd1 _0950_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_5_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0956__A1 _1100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0984_ _0971_/Y _1025_/A hold225/X _1071_/S vssd1 vssd1 vccd1 vccd1 _1554_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_13_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1605_ _1605_/CLK hold1/X _1387_/Y vssd1 vssd1 vccd1 vccd1 hold30/A sky130_fd_sc_hd__dfstp_1
X_1536_ _1556_/CLK _1536_/D _1318_/Y vssd1 vssd1 vccd1 vccd1 _1536_/Q sky130_fd_sc_hd__dfrtp_1
X_1467_ _1544_/CLK hold7/X _1249_/Y vssd1 vssd1 vccd1 vccd1 _1467_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1398_ _1409_/A vssd1 vssd1 vccd1 vccd1 _1398_/Y sky130_fd_sc_hd__inv_2
Xfanout128 _1416_/A vssd1 vssd1 vccd1 vccd1 _1402_/A sky130_fd_sc_hd__buf_4
Xfanout106 _1171_/S vssd1 vssd1 vccd1 vccd1 _1173_/S sky130_fd_sc_hd__buf_6
Xfanout117 _1007_/B vssd1 vssd1 vccd1 vccd1 _1100_/C sky130_fd_sc_hd__buf_4
XFILLER_0_54_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold115_A _0975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold193 _1434_/Q vssd1 vssd1 vccd1 vccd1 hold193/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 _1134_/X vssd1 vssd1 vccd1 vccd1 _1457_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold160 _1432_/Q vssd1 vssd1 vccd1 vccd1 hold160/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 hold180/X vssd1 vssd1 vccd1 vccd1 hold171/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1252_ _1415_/A vssd1 vssd1 vccd1 vccd1 _1252_/Y sky130_fd_sc_hd__inv_2
X_1321_ _1387_/A vssd1 vssd1 vccd1 vccd1 _1321_/Y sky130_fd_sc_hd__inv_2
X_1183_ _1183_/A _1183_/B vssd1 vssd1 vccd1 vccd1 _1183_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_46_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0967_ _1420_/Q _0967_/B _1418_/Q vssd1 vssd1 vccd1 vccd1 _0967_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_6_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0898_ _0897_/Y _0897_/A _0898_/S vssd1 vssd1 vccd1 vccd1 _1582_/D sky130_fd_sc_hd__mux2_1
X_1519_ _1634_/CLK _1519_/D _1301_/Y vssd1 vssd1 vccd1 vccd1 _1519_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0752_ hold2/X hold30/X _0752_/S vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__mux2_1
XFILLER_0_28_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0821_ _0817_/A _0816_/X _0820_/Y vssd1 vssd1 vccd1 vccd1 _0821_/X sky130_fd_sc_hd__o21a_1
XANTENNA__1024__B1 _1103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1235_ _1397_/A vssd1 vssd1 vccd1 vccd1 _1235_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1124__S _1135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1304_ _1417_/A vssd1 vssd1 vccd1 vccd1 _1304_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_29_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1166_ hold200/X hold218/X _1168_/S vssd1 vssd1 vccd1 vccd1 _1166_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1097_ input5/X input35/X input12/X input21/X _1007_/B _1100_/B vssd1 vssd1 vccd1
+ vccd1 _1098_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_19_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1006__B1 _1103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1020_ hold231/X _1059_/A2 _1103_/B _1019_/Y vssd1 vssd1 vccd1 vccd1 _1541_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_56_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0735_ _0741_/C _0882_/C vssd1 vssd1 vccd1 vccd1 _0735_/Y sky130_fd_sc_hd__nor2_1
X_0804_ _0837_/A _0837_/B _0804_/C _0804_/D vssd1 vssd1 vccd1 vccd1 _0813_/B sky130_fd_sc_hd__and4_1
XFILLER_0_21_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1119__S _1133_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1149_ hold263/X _1448_/Q _1168_/S vssd1 vssd1 vccd1 vccd1 _1149_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_46_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1218_ _1415_/A vssd1 vssd1 vccd1 vccd1 _1218_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_1_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold53 hold53/A vssd1 vssd1 vccd1 vccd1 hold53/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 hold64/A vssd1 vssd1 vccd1 vccd1 hold64/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 hold75/A vssd1 vssd1 vccd1 vccd1 hold75/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 hold86/A vssd1 vssd1 vccd1 vccd1 hold86/X sky130_fd_sc_hd__buf_2
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 hold97/A vssd1 vssd1 vccd1 vccd1 hold97/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1003_ hold6/X _1061_/A2 _1103_/B _1002_/X vssd1 vssd1 vccd1 vccd1 hold85/A sky130_fd_sc_hd__a22o_1
XFILLER_0_16_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0718_ _0826_/B vssd1 vssd1 vccd1 vccd1 _0776_/A sky130_fd_sc_hd__inv_2
XFILLER_0_12_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput98 _1461_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[5] sky130_fd_sc_hd__buf_12
Xoutput65 _1429_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[5] sky130_fd_sc_hd__buf_12
Xoutput54 _1448_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[24] sky130_fd_sc_hd__buf_12
Xoutput43 _1438_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[14] sky130_fd_sc_hd__buf_12
Xoutput76 _1470_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[14] sky130_fd_sc_hd__buf_12
Xoutput87 _1480_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[24] sky130_fd_sc_hd__buf_12
XFILLER_0_41_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1621_ _1625_/CLK _1621_/D _1403_/Y vssd1 vssd1 vccd1 vccd1 _1621_/Q sky130_fd_sc_hd__dfrtp_1
X_1552_ _1556_/CLK _1552_/D _1334_/Y vssd1 vssd1 vccd1 vccd1 _1552_/Q sky130_fd_sc_hd__dfrtp_1
X_1483_ _1582_/CLK _1483_/D _1265_/Y vssd1 vssd1 vccd1 vccd1 _1483_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1132__S _1135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold320 _0838_/X vssd1 vssd1 vccd1 vccd1 _1612_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 _1586_/Q vssd1 vssd1 vccd1 vccd1 hold375/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 _0808_/S vssd1 vssd1 vccd1 vccd1 _0810_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold342 _1623_/Q vssd1 vssd1 vccd1 vccd1 _0780_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold331 _1607_/Q vssd1 vssd1 vccd1 vccd1 hold331/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold386 _1419_/Q vssd1 vssd1 vccd1 vccd1 hold386/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold364 _1565_/Q vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0983_ _1100_/A _1007_/B _1007_/C vssd1 vssd1 vccd1 vccd1 _1025_/A sky130_fd_sc_hd__or3b_1
XANTENNA__1127__S _1133_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout107 _1135_/S vssd1 vssd1 vccd1 vccd1 _1133_/S sky130_fd_sc_hd__buf_6
Xfanout118 hold94/X vssd1 vssd1 vccd1 vccd1 _1007_/B sky130_fd_sc_hd__buf_4
Xfanout129 _1409_/A vssd1 vssd1 vccd1 vccd1 _1385_/A sky130_fd_sc_hd__buf_8
X_1604_ _1624_/CLK hold13/X _1386_/Y vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__dfrtp_1
X_1535_ _1556_/CLK _1535_/D _1317_/Y vssd1 vssd1 vccd1 vccd1 _1535_/Q sky130_fd_sc_hd__dfrtp_1
X_1397_ _1397_/A vssd1 vssd1 vccd1 vccd1 _1397_/Y sky130_fd_sc_hd__inv_2
X_1466_ _1547_/CLK _1466_/D _1248_/Y vssd1 vssd1 vccd1 vccd1 _1466_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1060__B2 _1031_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold194 _1163_/X vssd1 vssd1 vccd1 vccd1 _1434_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold150 _1026_/X vssd1 vssd1 vccd1 vccd1 _1538_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 _1522_/Q vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 _1165_/X vssd1 vssd1 vccd1 vccd1 _1432_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 _1127_/X vssd1 vssd1 vccd1 vccd1 _1464_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1320_ _1363_/A vssd1 vssd1 vccd1 vccd1 _1320_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1051__B2 _1031_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1251_ _1405_/A vssd1 vssd1 vccd1 vccd1 _1251_/Y sky130_fd_sc_hd__inv_2
X_1182_ _0847_/A _0784_/B _0852_/A _0836_/A _1101_/B vssd1 vssd1 vccd1 vccd1 _1182_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_46_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0897_ _0897_/A _0913_/A vssd1 vssd1 vccd1 vccd1 _0897_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_39_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1042__B2 _1059_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0966_ _1007_/B _0965_/Y _0966_/S vssd1 vssd1 vccd1 vccd1 _1561_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_49_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1518_ _1544_/CLK _1518_/D _1300_/Y vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__dfrtp_1
X_1449_ _1583_/CLK hold27/X _1231_/Y vssd1 vssd1 vccd1 vccd1 _1449_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_4_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1033__B2 _1030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1047__A2_N _1031_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0751_ _1583_/Q _0753_/D _1585_/Q _1584_/Q vssd1 vssd1 vccd1 vccd1 _0752_/S sky130_fd_sc_hd__and4bb_1
XFILLER_0_28_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0820_ _0865_/S _0820_/B vssd1 vssd1 vccd1 vccd1 _0820_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__1024__B2 _1023_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1303_ _1384_/A vssd1 vssd1 vccd1 vccd1 _1303_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_19_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1165_ hold131/X hold160/X _1168_/S vssd1 vssd1 vccd1 vccd1 _1165_/X sky130_fd_sc_hd__mux2_1
X_1234_ _1387_/A vssd1 vssd1 vccd1 vccd1 _1234_/Y sky130_fd_sc_hd__inv_2
X_1096_ _1095_/X hold60/X _1096_/S vssd1 vssd1 vccd1 vccd1 hold61/A sky130_fd_sc_hd__mux2_1
XANTENNA_fanout130_A _1416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0949_ hold86/X hold80/X _1100_/C vssd1 vssd1 vccd1 vccd1 _0955_/C sky130_fd_sc_hd__and3_1
XANTENNA__1006__B2 _1005_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0734_ _0917_/A _0734_/B vssd1 vssd1 vccd1 vccd1 _0882_/C sky130_fd_sc_hd__or2_2
X_0803_ _0803_/A _0817_/A _0822_/A _0803_/D vssd1 vssd1 vccd1 vccd1 _0804_/D sky130_fd_sc_hd__and4_1
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1135__S _1135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1148_ hold26/X _1449_/Q _1173_/S vssd1 vssd1 vccd1 vccd1 hold27/A sky130_fd_sc_hd__mux2_1
X_1217_ _1417_/A vssd1 vssd1 vccd1 vccd1 _1217_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_1_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1079_ input33/X input10/X input19/X input28/X _1100_/C _1100_/B vssd1 vssd1 vccd1
+ vccd1 _1080_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_30_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold54 hold54/A vssd1 vssd1 vccd1 vccd1 hold54/X sky130_fd_sc_hd__clkbuf_2
Xhold76 hold76/A vssd1 vssd1 vccd1 vccd1 hold76/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold43/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 hold87/A vssd1 vssd1 vccd1 vccd1 hold87/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 hold65/A vssd1 vssd1 vccd1 vccd1 hold65/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 hold98/A vssd1 vssd1 vccd1 vccd1 hold98/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold32/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1002_ hold81/X _1002_/B vssd1 vssd1 vccd1 vccd1 _1002_/X sky130_fd_sc_hd__and2_1
XFILLER_0_16_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0717_ _0886_/A vssd1 vssd1 vccd1 vccd1 _0717_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_57_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput55 _1449_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[25] sky130_fd_sc_hd__buf_12
Xoutput99 _1462_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[6] sky130_fd_sc_hd__buf_12
Xoutput88 _1481_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[25] sky130_fd_sc_hd__buf_12
Xoutput44 _1439_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[15] sky130_fd_sc_hd__buf_12
Xoutput77 _1471_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[15] sky130_fd_sc_hd__buf_12
Xoutput66 _1430_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[6] sky130_fd_sc_hd__buf_12
X_1620_ _1623_/CLK _1620_/D _1402_/Y vssd1 vssd1 vccd1 vccd1 _1620_/Q sky130_fd_sc_hd__dfrtp_1
X_1551_ _1634_/CLK hold83/X _1333_/Y vssd1 vssd1 vccd1 vccd1 hold76/A sky130_fd_sc_hd__dfrtp_1
X_1482_ _1600_/CLK _1482_/D _1264_/Y vssd1 vssd1 vccd1 vccd1 _1482_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_1_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold310 _0834_/X vssd1 vssd1 vccd1 vccd1 _1614_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold376 _1516_/Q vssd1 vssd1 vccd1 vccd1 hold376/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 _1609_/Q vssd1 vssd1 vccd1 vccd1 _0843_/A sky130_fd_sc_hd__buf_1
Xhold387 _1590_/Q vssd1 vssd1 vccd1 vccd1 hold84/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold354 _0810_/X vssd1 vssd1 vccd1 vccd1 _1622_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold343 _0808_/X vssd1 vssd1 vccd1 vccd1 _1623_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 _0856_/X vssd1 vssd1 vccd1 vccd1 _1607_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 _1603_/Q vssd1 vssd1 vccd1 vccd1 hold365/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0982_ _0971_/Y _1023_/A hold212/X _1061_/A2 vssd1 vssd1 vccd1 vccd1 _1555_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_13_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1534_ _1544_/CLK _1534_/D _1316_/Y vssd1 vssd1 vccd1 vccd1 _1534_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout108 _1129_/S vssd1 vssd1 vccd1 vccd1 _1135_/S sky130_fd_sc_hd__buf_6
X_1603_ _1624_/CLK hold15/X _1385_/Y vssd1 vssd1 vccd1 vccd1 _1603_/Q sky130_fd_sc_hd__dfrtp_1
Xfanout119 _1416_/A vssd1 vssd1 vccd1 vccd1 _1339_/A sky130_fd_sc_hd__buf_8
X_1465_ _1556_/CLK hold97/X _1247_/Y vssd1 vssd1 vccd1 vccd1 hold96/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1396_ _1397_/A vssd1 vssd1 vccd1 vccd1 _1396_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1143__S _1173_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold140 _0867_/X vssd1 vssd1 vccd1 vccd1 _1594_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 _1425_/Q vssd1 vssd1 vccd1 vccd1 hold151/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1060__A2 _1069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold162 hold388/X vssd1 vssd1 vccd1 vccd1 _1191_/B sky130_fd_sc_hd__clkbuf_2
Xhold184 _1429_/Q vssd1 vssd1 vccd1 vccd1 hold184/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 _1509_/Q vssd1 vssd1 vccd1 vccd1 hold195/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 _1564_/Q vssd1 vssd1 vccd1 vccd1 _0981_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_48_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1051__A2 _1069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1181_ hold336/X _1180_/X _1173_/S vssd1 vssd1 vccd1 vccd1 _1422_/D sky130_fd_sc_hd__a21bo_1
X_1250_ _1387_/A vssd1 vssd1 vccd1 vccd1 _1250_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_54_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0896_ _0896_/A _0933_/B _0905_/B _0896_/D vssd1 vssd1 vccd1 vccd1 _0898_/S sky130_fd_sc_hd__and4_1
XFILLER_0_42_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0965_ _1007_/B _1141_/B vssd1 vssd1 vccd1 vccd1 _0965_/Y sky130_fd_sc_hd__nor2_1
X_1448_ _1612_/CLK _1448_/D _1230_/Y vssd1 vssd1 vccd1 vccd1 _1448_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1517_ _1558_/CLK _1517_/D _1299_/Y vssd1 vssd1 vccd1 vccd1 hold34/A sky130_fd_sc_hd__dfrtp_1
X_1379_ _1402_/A vssd1 vssd1 vccd1 vccd1 _1379_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_52_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1033__A2 _1069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0750_ hold4/X hold30/X hold56/X vssd1 vssd1 vccd1 vccd1 hold57/A sky130_fd_sc_hd__mux2_1
XFILLER_0_24_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1024__A2 _1071_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1233_ _1404_/A vssd1 vssd1 vccd1 vccd1 _1233_/Y sky130_fd_sc_hd__inv_2
X_1302_ _1415_/A vssd1 vssd1 vccd1 vccd1 _1302_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_19_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1164_ hold286/X _1433_/Q _1168_/S vssd1 vssd1 vccd1 vccd1 _1164_/X sky130_fd_sc_hd__mux2_1
X_1095_ _1098_/A _1095_/B vssd1 vssd1 vccd1 vccd1 _1095_/X sky130_fd_sc_hd__and2_1
XFILLER_0_51_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0948_ _1100_/B _1007_/B vssd1 vssd1 vccd1 vccd1 _0963_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_15_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0879_ _0882_/A hold262/X hold56/X vssd1 vssd1 vccd1 vccd1 _1586_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_30_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1006__A2 _1059_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0802_ _0802_/A _0865_/S vssd1 vssd1 vccd1 vccd1 _0802_/Y sky130_fd_sc_hd__nor2_1
X_0733_ _0740_/A _0733_/B _0733_/C _0733_/D vssd1 vssd1 vccd1 vccd1 _0734_/B sky130_fd_sc_hd__or4_1
XANTENNA_clkbuf_leaf_3_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1216_ _1405_/A vssd1 vssd1 vccd1 vccd1 _1216_/Y sky130_fd_sc_hd__inv_2
X_1147_ hold72/X _1450_/Q _1173_/S vssd1 vssd1 vccd1 vccd1 hold73/A sky130_fd_sc_hd__mux2_1
XANTENNA__1046__A2_N _1031_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1151__S _1168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1078_ _1077_/X hold14/X _1099_/S vssd1 vssd1 vccd1 vccd1 _1496_/D sky130_fd_sc_hd__mux2_1
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 hold44/A vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 hold55/A vssd1 vssd1 vccd1 vccd1 hold55/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 hold77/A vssd1 vssd1 vccd1 vccd1 hold77/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 hold66/A vssd1 vssd1 vccd1 vccd1 hold66/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 hold88/A vssd1 vssd1 vccd1 vccd1 hold88/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 hold99/A vssd1 vssd1 vccd1 vccd1 hold99/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0986__B2 _1059_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1001_ _1100_/A _1100_/C hold84/X vssd1 vssd1 vccd1 vccd1 _1002_/B sky130_fd_sc_hd__and3b_1
XFILLER_0_29_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0716_ _0887_/B vssd1 vssd1 vccd1 vccd1 _0716_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1146__S _1168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0978__A1_N _0971_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput56 _1450_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[26] sky130_fd_sc_hd__buf_12
Xoutput89 _1482_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[26] sky130_fd_sc_hd__buf_12
Xoutput67 _1431_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[7] sky130_fd_sc_hd__buf_12
Xoutput78 _1472_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[16] sky130_fd_sc_hd__buf_12
Xoutput45 _1440_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[16] sky130_fd_sc_hd__buf_12
XFILLER_0_53_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0959__A1 _1100_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1550_ _1589_/CLK _1550_/D _1332_/Y vssd1 vssd1 vccd1 vccd1 hold52/A sky130_fd_sc_hd__dfrtp_1
X_1481_ _1544_/CLK _1481_/D _1263_/Y vssd1 vssd1 vccd1 vccd1 _1481_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold344 hold390/X vssd1 vssd1 vccd1 vccd1 _0919_/A sky130_fd_sc_hd__buf_1
Xhold300 _0734_/B vssd1 vssd1 vccd1 vccd1 _0736_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold322 _0844_/X vssd1 vssd1 vccd1 vccd1 _1609_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold311 _1621_/Q vssd1 vssd1 vccd1 vccd1 _0806_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold333 _1485_/Q vssd1 vssd1 vccd1 vccd1 hold333/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 _1567_/Q vssd1 vssd1 vccd1 vccd1 _0935_/S sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 _1531_/Q vssd1 vssd1 vccd1 vccd1 hold72/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 _1602_/Q vssd1 vssd1 vccd1 vccd1 hold366/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold388 _1593_/Q vssd1 vssd1 vccd1 vccd1 hold388/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1063__B1 _1027_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0981_ _0981_/A _1100_/C _1192_/B vssd1 vssd1 vccd1 vccd1 _1023_/A sky130_fd_sc_hd__or3b_1
XFILLER_0_13_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1602_ _1602_/CLK hold21/X _1384_/Y vssd1 vssd1 vccd1 vccd1 _1602_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1395_ _1397_/A vssd1 vssd1 vccd1 vccd1 _1395_/Y sky130_fd_sc_hd__inv_2
X_1464_ _1601_/CLK _1464_/D _1246_/Y vssd1 vssd1 vccd1 vccd1 _1464_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1533_ _1558_/CLK _1533_/D _1315_/Y vssd1 vssd1 vccd1 vccd1 hold98/A sky130_fd_sc_hd__dfrtp_1
Xfanout109 _1029_/X vssd1 vssd1 vccd1 vccd1 _1031_/C sky130_fd_sc_hd__buf_6
XFILLER_0_45_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold185 _1168_/X vssd1 vssd1 vccd1 vccd1 _1429_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 _0997_/X vssd1 vssd1 vccd1 vccd1 _1550_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold130 _1043_/X vssd1 vssd1 vccd1 vccd1 _1525_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 _1172_/X vssd1 vssd1 vccd1 vccd1 _1425_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 _1041_/X vssd1 vssd1 vccd1 vccd1 _1527_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 _1493_/Q vssd1 vssd1 vccd1 vccd1 hold141/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold196 _1059_/X vssd1 vssd1 vccd1 vccd1 _1509_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_21_clk clkbuf_1_1__f_clk/X vssd1 vssd1 vccd1 vccd1 _1600_/CLK sky130_fd_sc_hd__clkbuf_16
X_1180_ _1180_/A _1180_/B _1183_/B vssd1 vssd1 vccd1 vccd1 _1180_/X sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_12_clk clkbuf_1_1__f_clk/X vssd1 vssd1 vccd1 vccd1 _1612_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_42_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0964_ _1100_/B _0963_/X _0966_/S vssd1 vssd1 vccd1 vccd1 _1562_/D sky130_fd_sc_hd__mux2_1
X_0895_ _0896_/A _0905_/B _0896_/D vssd1 vssd1 vccd1 vccd1 _0895_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_42_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1516_ _1589_/CLK _1516_/D _1298_/Y vssd1 vssd1 vccd1 vccd1 _1516_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1154__S _1173_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1447_ _1615_/CLK _1447_/D _1229_/Y vssd1 vssd1 vccd1 vccd1 _1447_/Q sky130_fd_sc_hd__dfrtp_1
X_1378_ _1402_/A vssd1 vssd1 vccd1 vccd1 _1378_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_10_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1018__B1 _1103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1064__S _1071_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1009__B1 _1103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1232_ _1417_/A vssd1 vssd1 vccd1 vccd1 _1232_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_1_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _1634_/CLK sky130_fd_sc_hd__clkbuf_16
X_1301_ _1415_/A vssd1 vssd1 vccd1 vccd1 _1301_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_19_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1163_ hold126/X hold193/X _1168_/S vssd1 vssd1 vccd1 vccd1 _1163_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_35_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1094_ input16/X input36/X input13/X input22/X _1100_/C _1100_/B vssd1 vssd1 vccd1
+ vccd1 _1095_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_51_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1149__S _1168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0947_ _1179_/A _0947_/B _0947_/C vssd1 vssd1 vccd1 vccd1 _0966_/S sky130_fd_sc_hd__and3b_2
XFILLER_0_42_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0878_ _0933_/B hold55/X _0880_/B vssd1 vssd1 vccd1 vccd1 _0878_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_33_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0801_ _0826_/B _0801_/B vssd1 vssd1 vccd1 vccd1 _0836_/A sky130_fd_sc_hd__or2_2
X_0732_ _0914_/S _0912_/A _0919_/A _1573_/Q vssd1 vssd1 vccd1 vccd1 _0733_/D sky130_fd_sc_hd__or4b_1
XFILLER_0_12_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1146_ hold58/X hold78/X _1168_/S vssd1 vssd1 vccd1 vccd1 hold79/A sky130_fd_sc_hd__mux2_1
X_1215_ _1385_/A vssd1 vssd1 vccd1 vccd1 _1215_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1077_ _1098_/A _1077_/B vssd1 vssd1 vccd1 vccd1 _1077_/X sky130_fd_sc_hd__and2_1
XFILLER_0_30_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 hold56/A vssd1 vssd1 vccd1 vccd1 hold56/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 hold78/A vssd1 vssd1 vccd1 vccd1 hold78/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 hold67/A vssd1 vssd1 vccd1 vccd1 hold67/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 hold89/A vssd1 vssd1 vccd1 vccd1 hold89/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1000_ hold220/X _1071_/S _1103_/B _0999_/X vssd1 vssd1 vccd1 vccd1 _1549_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0715_ _0892_/B vssd1 vssd1 vccd1 vccd1 _0910_/A sky130_fd_sc_hd__inv_2
XFILLER_0_57_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1129_ hold110/X hold204/X _1129_/S vssd1 vssd1 vccd1 vccd1 _1129_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1162__S _1173_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput57 hold78/A vssd1 vssd1 vccd1 vccd1 wb_adr_o[27] sky130_fd_sc_hd__buf_12
XFILLER_0_43_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput46 _1441_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[17] sky130_fd_sc_hd__buf_12
Xoutput79 _1473_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[17] sky130_fd_sc_hd__buf_12
Xoutput68 _1432_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[8] sky130_fd_sc_hd__buf_12
XANTENNA_clkbuf_leaf_2_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0959__A2 _1100_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1045__A2_N _1031_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1480_ _1605_/CLK _1480_/D _1262_/Y vssd1 vssd1 vccd1 vccd1 _1480_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1011__A hold81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold301 _1579_/Q vssd1 vssd1 vccd1 vccd1 _0905_/A sky130_fd_sc_hd__buf_1
Xhold334 _1577_/Q vssd1 vssd1 vccd1 vccd1 _0892_/B sky130_fd_sc_hd__buf_1
Xhold345 _0906_/B vssd1 vssd1 vccd1 vccd1 hold345/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 _1573_/Q vssd1 vssd1 vccd1 vccd1 _0923_/S sky130_fd_sc_hd__buf_1
XFILLER_0_40_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold378 _1589_/Q vssd1 vssd1 vccd1 vccd1 hold378/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 _1594_/Q vssd1 vssd1 vccd1 vccd1 hold367/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 _1616_/Q vssd1 vssd1 vccd1 vccd1 _0803_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold312 _0773_/X vssd1 vssd1 vccd1 vccd1 _0774_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1157__S _1168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold389 _1563_/Q vssd1 vssd1 vccd1 vccd1 hold86/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1063__B2 _1031_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1067__S _1071_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0980_ _0971_/Y _1021_/A hold22/X _1069_/S vssd1 vssd1 vccd1 vccd1 hold95/A sky130_fd_sc_hd__a2bb2o_1
XANTENNA__1054__A1 hold286/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1054__B2 _1031_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1532_ _1548_/CLK hold59/X _1314_/Y vssd1 vssd1 vccd1 vccd1 hold58/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1601_ _1601_/CLK hold63/X _1383_/Y vssd1 vssd1 vccd1 vccd1 hold62/A sky130_fd_sc_hd__dfrtp_1
X_1463_ _1582_/CLK _1463_/D _1245_/Y vssd1 vssd1 vccd1 vccd1 _1463_/Q sky130_fd_sc_hd__dfrtp_1
X_1394_ _1397_/A vssd1 vssd1 vccd1 vccd1 _1394_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_38_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold175 _1560_/Q vssd1 vssd1 vccd1 vccd1 hold175/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 hold375/X vssd1 vssd1 vccd1 vccd1 _0882_/A sky130_fd_sc_hd__buf_1
Xhold153 _1489_/Q vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 _1513_/Q vssd1 vssd1 vccd1 vccd1 hold131/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 _1595_/Q vssd1 vssd1 vccd1 vccd1 _1140_/A sky130_fd_sc_hd__buf_2
XFILLER_0_0_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold186 _1466_/Q vssd1 vssd1 vccd1 vccd1 hold186/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 _1087_/X vssd1 vssd1 vccd1 vccd1 _1493_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 _1496_/Q vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1036__B2 _1030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0894_ _0905_/B _0896_/D vssd1 vssd1 vccd1 vccd1 _0894_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_39_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0963_ _0963_/A _0963_/B _0963_/C vssd1 vssd1 vccd1 vccd1 _0963_/X sky130_fd_sc_hd__and3_1
XFILLER_0_57_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1515_ _1544_/CLK _1515_/D _1297_/Y vssd1 vssd1 vccd1 vccd1 _1515_/Q sky130_fd_sc_hd__dfrtp_1
X_1377_ _1410_/A vssd1 vssd1 vccd1 vccd1 _1377_/Y sky130_fd_sc_hd__inv_2
X_1446_ _1547_/CLK hold71/X _1228_/Y vssd1 vssd1 vccd1 vccd1 _1446_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1170__S _1173_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1300_ _1405_/A vssd1 vssd1 vccd1 vccd1 _1300_/Y sky130_fd_sc_hd__inv_2
X_1231_ _1363_/A vssd1 vssd1 vccd1 vccd1 _1231_/Y sky130_fd_sc_hd__inv_2
X_1162_ hold265/X _1435_/Q _1173_/S vssd1 vssd1 vccd1 vccd1 _1162_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_35_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1093_ _1092_/X hold135/X _1099_/S vssd1 vssd1 vccd1 vccd1 _1491_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_19_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0877_ _0917_/A _0741_/C hold345/X _0919_/B vssd1 vssd1 vccd1 vccd1 _0880_/B sky130_fd_sc_hd__o31a_1
XFILLER_0_30_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0946_ _1141_/A _1140_/A _0946_/C vssd1 vssd1 vccd1 vccd1 _0947_/C sky130_fd_sc_hd__or3_1
X_1429_ _1612_/CLK _1429_/D _1211_/Y vssd1 vssd1 vccd1 vccd1 _1429_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1165__S _1168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout109_A _1029_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0731_ _0889_/C _1571_/Q _0731_/C _1568_/Q vssd1 vssd1 vccd1 vccd1 _0731_/X sky130_fd_sc_hd__or4_1
X_0800_ _1606_/Q _0801_/B vssd1 vssd1 vccd1 vccd1 _0865_/S sky130_fd_sc_hd__nor2_4
XFILLER_0_21_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1214_ _1409_/A vssd1 vssd1 vccd1 vccd1 _1214_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_1_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1145_ hold98/X _1452_/Q _1173_/S vssd1 vssd1 vccd1 vccd1 hold99/A sky130_fd_sc_hd__mux2_1
XFILLER_0_1_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1076_ input34/X input11/X input20/X input29/X _1100_/C _1100_/B vssd1 vssd1 vccd1
+ vccd1 _1077_/B sky130_fd_sc_hd__mux4_1
X_0929_ _0717_/Y _0885_/Y _0928_/X vssd1 vssd1 vccd1 vccd1 _0929_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 hold68/A vssd1 vssd1 vccd1 vccd1 hold68/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 hold79/A vssd1 vssd1 vccd1 vccd1 hold79/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 hold57/A vssd1 vssd1 vccd1 vccd1 hold57/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold173_A _1564_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 hold35/A vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0714_ _0739_/A vssd1 vssd1 vccd1 vccd1 _0897_/A sky130_fd_sc_hd__inv_2
XFILLER_0_4_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1128_ hold259/X _1463_/Q _1129_/S vssd1 vssd1 vccd1 vccd1 _1128_/X sky130_fd_sc_hd__mux2_1
X_1059_ hold195/X _1059_/A2 _1019_/Y hold165/X vssd1 vssd1 vccd1 vccd1 _1059_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput47 _1442_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[18] sky130_fd_sc_hd__buf_12
Xoutput58 _1452_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[28] sky130_fd_sc_hd__buf_12
XFILLER_0_9_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput69 _1433_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[9] sky130_fd_sc_hd__buf_12
XFILLER_0_34_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold335 _0911_/Y vssd1 vssd1 vccd1 vccd1 _1577_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold302 _0907_/X vssd1 vssd1 vccd1 vccd1 _1579_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 _0923_/X vssd1 vssd1 vccd1 vccd1 _1573_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold357 _0824_/X vssd1 vssd1 vccd1 vccd1 _0825_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold368 _1598_/Q vssd1 vssd1 vccd1 vccd1 hold368/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold379 _1587_/Q vssd1 vssd1 vccd1 vccd1 hold379/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold313 _0784_/B vssd1 vssd1 vccd1 vccd1 hold313/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold346 _1418_/Q vssd1 vssd1 vccd1 vccd1 hold346/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1173__S _1173_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1063__A2 _1069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1054__A2 _1069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1462_ _1544_/CLK _1462_/D _1244_/Y vssd1 vssd1 vccd1 vccd1 _1462_/Q sky130_fd_sc_hd__dfrtp_4
X_1531_ _1548_/CLK _1531_/D _1313_/Y vssd1 vssd1 vccd1 vccd1 _1531_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1600_ _1600_/CLK _1600_/D _1382_/Y vssd1 vssd1 vccd1 vccd1 _1600_/Q sky130_fd_sc_hd__dfrtp_1
X_1393_ _1397_/A vssd1 vssd1 vccd1 vccd1 _1393_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_57_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1168__S _1168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold110 _1543_/Q vssd1 vssd1 vccd1 vccd1 hold110/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 _1112_/X vssd1 vssd1 vccd1 vccd1 _1479_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 _1542_/Q vssd1 vssd1 vccd1 vccd1 hold154/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 hold373/X vssd1 vssd1 vccd1 vccd1 _1007_/C sky130_fd_sc_hd__clkbuf_2
Xhold198 _0874_/S vssd1 vssd1 vccd1 vccd1 _1595_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 hold374/X vssd1 vssd1 vccd1 vccd1 _0989_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_1_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold132 _1055_/X vssd1 vssd1 vccd1 vccd1 _1513_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 _1125_/X vssd1 vssd1 vccd1 vccd1 _1466_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 _1029_/X vssd1 vssd1 vccd1 vccd1 hold165/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1044__A2_N _1031_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0893_ _0893_/A _0905_/A vssd1 vssd1 vccd1 vccd1 _0896_/D sky130_fd_sc_hd__and2_1
XFILLER_0_42_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0962_ _1100_/B _1007_/B vssd1 vssd1 vccd1 vccd1 _0963_/C sky130_fd_sc_hd__or2_1
XFILLER_0_49_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1017__A _1017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1445_ _1547_/CLK hold43/X _1227_/Y vssd1 vssd1 vccd1 vccd1 _1445_/Q sky130_fd_sc_hd__dfrtp_1
X_1514_ _1556_/CLK _1514_/D _1296_/Y vssd1 vssd1 vccd1 vccd1 _1514_/Q sky130_fd_sc_hd__dfrtp_1
X_1376_ _1417_/A vssd1 vssd1 vccd1 vccd1 _1376_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1018__A2 _1059_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0976__A1_N _0971_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1009__A2 _1069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1230_ _1397_/A vssd1 vssd1 vccd1 vccd1 _1230_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_35_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1092_ _1098_/A _1092_/B vssd1 vssd1 vccd1 vccd1 _1092_/X sky130_fd_sc_hd__and2_1
X_1161_ hold34/X _1436_/Q _1173_/S vssd1 vssd1 vccd1 vccd1 hold35/A sky130_fd_sc_hd__mux2_1
XFILLER_0_19_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0876_ _0919_/B vssd1 vssd1 vccd1 vccd1 _0913_/A sky130_fd_sc_hd__inv_2
XFILLER_0_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0945_ _1101_/C _1185_/A _1185_/B _0945_/D vssd1 vssd1 vccd1 vccd1 _0947_/B sky130_fd_sc_hd__or4_1
X_1428_ _1612_/CLK _1428_/D _1210_/Y vssd1 vssd1 vccd1 vccd1 _1428_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1359_ _1364_/A vssd1 vssd1 vccd1 vccd1 _1359_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_33_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0730_ _0739_/A _1581_/Q _1569_/Q _1567_/Q vssd1 vssd1 vccd1 vccd1 _0730_/X sky130_fd_sc_hd__or4bb_1
X_1213_ _1385_/A vssd1 vssd1 vccd1 vccd1 _1213_/Y sky130_fd_sc_hd__inv_2
X_1144_ hold253/X _1453_/Q _1168_/S vssd1 vssd1 vccd1 vccd1 _1144_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1075_ _1100_/A hold86/X _1101_/C vssd1 vssd1 vccd1 vccd1 _1098_/A sky130_fd_sc_hd__nor3b_4
XFILLER_0_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout121_A _1416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0928_ _0886_/A _0925_/A _0915_/C _0917_/A vssd1 vssd1 vccd1 vccd1 _0928_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_30_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0859_ hold366/X hold20/X _0865_/S vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__mux2_1
Xhold47 hold47/A vssd1 vssd1 vccd1 vccd1 hold47/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 hold69/A vssd1 vssd1 vccd1 vccd1 hold69/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 hold58/A vssd1 vssd1 vccd1 vccd1 hold58/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0713_ _0884_/S vssd1 vssd1 vccd1 vccd1 _0764_/B sky130_fd_sc_hd__inv_2
XFILLER_0_12_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1058_ hold158/X _1061_/A2 _1017_/Y _1029_/X vssd1 vssd1 vccd1 vccd1 _1058_/X sky130_fd_sc_hd__a22o_1
X_1127_ hold171/X _1464_/Q _1133_/S vssd1 vssd1 vccd1 vccd1 _1127_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_35_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput37 _1607_/Q vssd1 vssd1 vccd1 vccd1 o_uart_tx sky130_fd_sc_hd__buf_12
Xoutput59 _1453_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[29] sky130_fd_sc_hd__buf_12
Xoutput48 _1443_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[19] sky130_fd_sc_hd__buf_12
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1066__A0 _0995_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1057__B1 _1015_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold303 _1569_/Q vssd1 vssd1 vccd1 vccd1 _0886_/B sky130_fd_sc_hd__buf_1
Xhold347 _1571_/Q vssd1 vssd1 vccd1 vccd1 _0887_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold358 _0825_/X vssd1 vssd1 vccd1 vccd1 _1616_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 _1596_/Q vssd1 vssd1 vccd1 vccd1 hold369/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold336 _1636_/A vssd1 vssd1 vccd1 vccd1 hold336/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold325 _1486_/Q vssd1 vssd1 vccd1 vccd1 hold325/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold314 _0787_/X vssd1 vssd1 vccd1 vccd1 _1627_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_24_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _1562_/CLK sky130_fd_sc_hd__clkbuf_16
X_1461_ _1612_/CLK _1461_/D _1243_/Y vssd1 vssd1 vccd1 vccd1 _1461_/Q sky130_fd_sc_hd__dfrtp_1
X_1530_ _1586_/CLK _1530_/D _1312_/Y vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1392_ _1404_/A vssd1 vssd1 vccd1 vccd1 _1392_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_22_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_15_clk clkbuf_1_1__f_clk/X vssd1 vssd1 vccd1 vccd1 _1598_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold111 _1016_/X vssd1 vssd1 vccd1 vccd1 _1543_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 _1007_/X vssd1 vssd1 vccd1 vccd1 _1008_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 _1456_/Q vssd1 vssd1 vccd1 vccd1 hold133/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold100 _1520_/Q vssd1 vssd1 vccd1 vccd1 hold100/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold144 _0990_/B vssd1 vssd1 vccd1 vccd1 hold144/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold155 _1018_/X vssd1 vssd1 vccd1 vccd1 _1542_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 _0870_/X vssd1 vssd1 vccd1 vccd1 _1591_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 hold386/X vssd1 vssd1 vccd1 vccd1 _0967_/B sky130_fd_sc_hd__buf_2
Xhold166 _1060_/X vssd1 vssd1 vccd1 vccd1 _1508_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 _1471_/Q vssd1 vssd1 vccd1 vccd1 hold188/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0962__A _1100_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0961_ hold86/X _0960_/X _0966_/S vssd1 vssd1 vccd1 vccd1 _1563_/D sky130_fd_sc_hd__mux2_1
X_0892_ _0892_/A _0892_/B _0910_/C vssd1 vssd1 vccd1 vccd1 _0905_/B sky130_fd_sc_hd__and3_2
XFILLER_0_54_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1017__B _1027_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1444_ _1612_/CLK hold51/X _1226_/Y vssd1 vssd1 vccd1 vccd1 _1444_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_4_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _1635_/CLK sky130_fd_sc_hd__clkbuf_16
X_1375_ _1415_/A vssd1 vssd1 vccd1 vccd1 _1375_/Y sky130_fd_sc_hd__inv_2
X_1513_ _1627_/CLK _1513_/D _1295_/Y vssd1 vssd1 vccd1 vccd1 _1513_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1193__A2 _1191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1160_ hold46/X _1437_/Q _1168_/S vssd1 vssd1 vccd1 vccd1 hold47/A sky130_fd_sc_hd__mux2_1
X_1091_ input27/X input6/X input14/X input23/X _1007_/B _1100_/B vssd1 vssd1 vccd1
+ vccd1 _1092_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_35_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_0_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0944_ _1141_/A _1180_/A vssd1 vssd1 vccd1 vccd1 _0945_/D sky130_fd_sc_hd__nor2_1
X_0875_ input1/X _0917_/A vssd1 vssd1 vccd1 vccd1 _0919_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_2_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1358_ _1364_/A vssd1 vssd1 vccd1 vccd1 _1358_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1043__A2_N _1031_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1427_ _1505_/CLK hold89/X _1209_/Y vssd1 vssd1 vccd1 vccd1 _1427_/Q sky130_fd_sc_hd__dfrtp_1
X_1289_ _1324_/A vssd1 vssd1 vccd1 vccd1 _1289_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_33_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1212_ _1385_/A vssd1 vssd1 vccd1 vccd1 _1212_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_1_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1143_ hold236/X hold250/X _1173_/S vssd1 vssd1 vccd1 vccd1 _1143_/X sky130_fd_sc_hd__mux2_1
X_1074_ _1101_/C hold107/X _1183_/A _1073_/Y vssd1 vssd1 vccd1 vccd1 _1096_/S sky130_fd_sc_hd__a211o_1
X_0927_ _0716_/Y _0925_/Y _0925_/B _0915_/C vssd1 vssd1 vccd1 vccd1 _1571_/D sky130_fd_sc_hd__a2bb2o_1
XANTENNA__1030__B _1100_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0858_ hold365/X hold14/X _0865_/S vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__mux2_1
X_0789_ _0789_/A _0851_/S vssd1 vssd1 vccd1 vccd1 _0789_/X sky130_fd_sc_hd__or2_1
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 hold59/A vssd1 vssd1 vccd1 vccd1 hold59/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 hold48/A vssd1 vssd1 vccd1 vccd1 hold48/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0712_ _0764_/A vssd1 vssd1 vccd1 vccd1 _0754_/A sky130_fd_sc_hd__inv_2
XFILLER_0_12_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1025__B _1027_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1126_ hold90/X hold96/X _1133_/S vssd1 vssd1 vccd1 vccd1 hold97/A sky130_fd_sc_hd__mux2_1
X_1057_ hold36/X _1059_/A2 _1015_/Y _1031_/C vssd1 vssd1 vccd1 vccd1 _1511_/D sky130_fd_sc_hd__a22o_1
Xoutput49 _1425_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[1] sky130_fd_sc_hd__buf_12
Xoutput38 _1424_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[0] sky130_fd_sc_hd__buf_12
XFILLER_0_11_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0965__A _1007_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1057__B2 _1031_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold315 _1581_/Q vssd1 vssd1 vccd1 vccd1 _0896_/A sky130_fd_sc_hd__buf_1
Xhold326 _1483_/Q vssd1 vssd1 vccd1 vccd1 hold326/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold304 _0931_/X vssd1 vssd1 vccd1 vccd1 _1569_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold348 _1570_/Q vssd1 vssd1 vccd1 vccd1 _0731_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 _1617_/Q vssd1 vssd1 vccd1 vccd1 _0822_/A sky130_fd_sc_hd__buf_1
Xhold359 _1606_/Q vssd1 vssd1 vccd1 vccd1 _0826_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_7_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1109_ _1192_/B hold305/X _1133_/S vssd1 vssd1 vccd1 vccd1 _1482_/D sky130_fd_sc_hd__mux2_1
XANTENNA__1048__B2 _1031_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1039__B2 _1030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1460_ _1612_/CLK _1460_/D _1242_/Y vssd1 vssd1 vccd1 vccd1 _1460_/Q sky130_fd_sc_hd__dfrtp_1
X_1391_ _1404_/A vssd1 vssd1 vccd1 vccd1 _1391_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_54_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0957__A_N _1100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold167 _1461_/Q vssd1 vssd1 vccd1 vccd1 hold167/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 _1038_/X vssd1 vssd1 vccd1 vccd1 _1530_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 _1135_/X vssd1 vssd1 vccd1 vccd1 _1456_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 _1537_/Q vssd1 vssd1 vccd1 vccd1 hold112/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold101 _1158_/X vssd1 vssd1 vccd1 vccd1 _1439_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 _1547_/Q vssd1 vssd1 vccd1 vccd1 hold156/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 _1048_/X vssd1 vssd1 vccd1 vccd1 _1520_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1589_ _1589_/CLK hold17/X _1371_/Y vssd1 vssd1 vccd1 vccd1 _1589_/Q sky130_fd_sc_hd__dfrtp_1
Xhold178 _0967_/Y vssd1 vssd1 vccd1 vccd1 _1073_/B sky130_fd_sc_hd__buf_1
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold189 _1120_/X vssd1 vssd1 vccd1 vccd1 _1471_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1177__B1_N _1135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0962__B _1007_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0960_ _0955_/C _0963_/B _0960_/C _0960_/D vssd1 vssd1 vccd1 vccd1 _0960_/X sky130_fd_sc_hd__and4b_1
X_0891_ _0892_/B _0910_/C vssd1 vssd1 vccd1 vccd1 _0891_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_40_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1512_ _1601_/CLK _1512_/D _1294_/Y vssd1 vssd1 vccd1 vccd1 _1512_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1443_ _1583_/CLK hold29/X _1225_/Y vssd1 vssd1 vccd1 vccd1 _1443_/Q sky130_fd_sc_hd__dfrtp_1
X_1374_ _1415_/A vssd1 vssd1 vccd1 vccd1 _1374_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_14_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1178__A0 _1031_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1090_ _1089_/X hold214/X _1099_/S vssd1 vssd1 vccd1 vccd1 _1090_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0973__A _1100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0874_ hold370/X hold40/X _0874_/S vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__mux2_1
XFILLER_0_27_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0943_ _1141_/A _0967_/B _1180_/A vssd1 vssd1 vccd1 vccd1 _1185_/B sky130_fd_sc_hd__and3b_1
XFILLER_0_50_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1357_ _1364_/A vssd1 vssd1 vccd1 vccd1 _1357_/Y sky130_fd_sc_hd__inv_2
X_1426_ _1612_/CLK hold69/X _1208_/Y vssd1 vssd1 vccd1 vccd1 _1426_/Q sky130_fd_sc_hd__dfrtp_2
X_1288_ _1417_/A vssd1 vssd1 vccd1 vccd1 _1288_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_33_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1211_ _1397_/A vssd1 vssd1 vccd1 vccd1 _1211_/Y sky130_fd_sc_hd__inv_2
X_1142_ hold234/X _1455_/Q _1173_/S vssd1 vssd1 vccd1 vccd1 _1142_/X sky130_fd_sc_hd__mux2_1
X_1073_ _1101_/C _1073_/B vssd1 vssd1 vccd1 vccd1 _1073_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_1_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0926_ _0917_/A _0917_/B _0925_/Y _0889_/C vssd1 vssd1 vccd1 vccd1 _0926_/X sky130_fd_sc_hd__o22a_1
XANTENNA__1030__C _1031_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0857_ hold12/X _0865_/S vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__or2_1
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1409_ _1409_/A vssd1 vssd1 vccd1 vccd1 _1409_/Y sky130_fd_sc_hd__inv_2
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout107_A _1135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0788_ _0768_/B _0784_/X _0785_/X _0850_/A vssd1 vssd1 vccd1 vccd1 _0788_/X sky130_fd_sc_hd__a22o_1
Xhold49 hold49/A vssd1 vssd1 vccd1 vccd1 hold49/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0711_ hold54/X vssd1 vssd1 vccd1 vccd1 _0753_/A sky130_fd_sc_hd__inv_2
XANTENNA__1042__A2_N _1031_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1125_ hold156/X hold186/X _1133_/S vssd1 vssd1 vccd1 vccd1 _1125_/X sky130_fd_sc_hd__mux2_1
X_1056_ hold200/X _1059_/A2 _1013_/Y _1031_/C vssd1 vssd1 vccd1 vccd1 _1056_/X sky130_fd_sc_hd__a22o_1
Xoutput39 _1434_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[10] sky130_fd_sc_hd__buf_12
X_0909_ _1566_/Q _0905_/B _0908_/Y _0892_/A vssd1 vssd1 vccd1 vccd1 _0909_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_43_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0949__C _1100_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0974__A1_N _0971_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1057__A2 _1059_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold316 _0901_/X vssd1 vssd1 vccd1 vccd1 _1581_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 _0731_/X vssd1 vssd1 vccd1 vccd1 _0733_/C sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold338 _0822_/Y vssd1 vssd1 vccd1 vccd1 hold338/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold327 _1484_/Q vssd1 vssd1 vccd1 vccd1 hold327/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold305 _1482_/Q vssd1 vssd1 vccd1 vccd1 hold305/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1108_ hold84/X hold326/X _1135_/S vssd1 vssd1 vccd1 vccd1 _1483_/D sky130_fd_sc_hd__mux2_1
X_1039_ hold263/X _1061_/A2 _1011_/B _1030_/X vssd1 vssd1 vccd1 vccd1 _1529_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1048__A2 _1069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1390_ _1397_/A vssd1 vssd1 vccd1 vccd1 _1390_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_54_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold168 _1130_/X vssd1 vssd1 vccd1 vccd1 _1461_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 _1028_/X vssd1 vssd1 vccd1 vccd1 _1537_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1588_ _1631_/CLK _1588_/D _1370_/Y vssd1 vssd1 vccd1 vccd1 _1588_/Q sky130_fd_sc_hd__dfrtp_1
Xhold146 _1491_/Q vssd1 vssd1 vccd1 vccd1 hold146/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 hold146/X vssd1 vssd1 vccd1 vccd1 hold135/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold102 _1424_/Q vssd1 vssd1 vccd1 vccd1 hold102/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 _1006_/X vssd1 vssd1 vccd1 vccd1 _1547_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold179 _1035_/X vssd1 vssd1 vccd1 vccd1 _1533_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 _1600_/Q vssd1 vssd1 vccd1 vccd1 hold124/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0890_ _0914_/S _0912_/A _0915_/C _0915_/D vssd1 vssd1 vccd1 vccd1 _0910_/C sky130_fd_sc_hd__and4_1
XFILLER_0_42_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1442_ _1625_/CLK _1442_/D _1224_/Y vssd1 vssd1 vccd1 vccd1 _1442_/Q sky130_fd_sc_hd__dfrtp_1
X_1511_ _1624_/CLK _1511_/D _1293_/Y vssd1 vssd1 vccd1 vccd1 hold36/A sky130_fd_sc_hd__dfrtp_1
X_1373_ _1410_/A vssd1 vssd1 vccd1 vccd1 _1373_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_18_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0957__C _1100_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0973__B _1100_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0873_ _1007_/C hold210/X _0874_/S vssd1 vssd1 vccd1 vccd1 _0873_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0942_ _0967_/B _1180_/A _1141_/A vssd1 vssd1 vccd1 vccd1 _1185_/A sky130_fd_sc_hd__and3b_1
XFILLER_0_50_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1425_ _1586_/CLK _1425_/D _1207_/Y vssd1 vssd1 vccd1 vccd1 _1425_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1356_ _1364_/A vssd1 vssd1 vccd1 vccd1 _1356_/Y sky130_fd_sc_hd__inv_2
X_1287_ _1339_/A vssd1 vssd1 vccd1 vccd1 _1287_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_25_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0983__C_N _1007_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1020__B1 _1103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1210_ _1397_/A vssd1 vssd1 vccd1 vccd1 _1210_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_46_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1072_ _1140_/A _1073_/B vssd1 vssd1 vccd1 vccd1 _1183_/A sky130_fd_sc_hd__and2b_1
X_1141_ _1141_/A _1141_/B _1141_/C _1141_/D vssd1 vssd1 vccd1 vccd1 _1171_/S sky130_fd_sc_hd__or4_4
XFILLER_0_55_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0925_ _0925_/A _0925_/B vssd1 vssd1 vccd1 vccd1 _0925_/Y sky130_fd_sc_hd__nor2_1
X_0856_ hold331/X _0783_/X _0855_/X hold313/X vssd1 vssd1 vccd1 vccd1 _0856_/X sky130_fd_sc_hd__a22o_1
X_0787_ _0847_/A _0785_/X _0786_/Y hold313/X vssd1 vssd1 vccd1 vccd1 _0787_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_11_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__dlygate4sd3_1
X_1408_ _1409_/A vssd1 vssd1 vccd1 vccd1 _1408_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_38_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1339_ _1339_/A vssd1 vssd1 vccd1 vccd1 _1339_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0979__A _1100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0710_ _0989_/C vssd1 vssd1 vccd1 vccd1 _1191_/A sky130_fd_sc_hd__inv_2
XFILLER_0_12_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1124_ hold6/X _1467_/Q _1135_/S vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__mux2_1
X_1055_ hold131/X _1059_/A2 _1011_/X _1031_/C vssd1 vssd1 vccd1 vccd1 _1055_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_22_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0908_ _0933_/B _0891_/Y _0925_/A vssd1 vssd1 vccd1 vccd1 _0908_/Y sky130_fd_sc_hd__a21oi_1
X_0839_ _1610_/Q _1609_/Q _1608_/Q _0795_/A vssd1 vssd1 vccd1 vccd1 _0839_/X sky130_fd_sc_hd__a31o_1
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_27_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _1505_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_43_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0981__B _1100_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold328 _1568_/Q vssd1 vssd1 vccd1 vccd1 _0886_/C sky130_fd_sc_hd__buf_1
XFILLER_0_40_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold339 _0823_/Y vssd1 vssd1 vccd1 vccd1 _1617_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold306 _1480_/Q vssd1 vssd1 vccd1 vccd1 hold306/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold317 _1624_/Q vssd1 vssd1 vccd1 vccd1 _0851_/S sky130_fd_sc_hd__buf_2
X_1038_ hold26/X _1071_/S _1008_/B _1030_/X vssd1 vssd1 vccd1 vccd1 _1038_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_18_clk clkbuf_1_1__f_clk/X vssd1 vssd1 vccd1 vccd1 _1624_/CLK sky130_fd_sc_hd__clkbuf_16
X_1107_ _1192_/D hold327/X _1133_/S vssd1 vssd1 vccd1 vccd1 _1484_/D sky130_fd_sc_hd__mux2_1
XANTENNA__1041__A2_N _1031_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_7_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _1582_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold158 _1510_/Q vssd1 vssd1 vccd1 vccd1 hold158/X sky130_fd_sc_hd__dlygate4sd3_1
X_1587_ _1631_/CLK hold41/X _1369_/Y vssd1 vssd1 vccd1 vccd1 _1587_/Q sky130_fd_sc_hd__dfrtp_1
Xhold136 _0863_/X vssd1 vssd1 vccd1 vccd1 _1598_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold169 _1458_/Q vssd1 vssd1 vccd1 vccd1 hold169/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold103 _1173_/X vssd1 vssd1 vccd1 vccd1 _1424_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 _1552_/Q vssd1 vssd1 vccd1 vccd1 hold147/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold125 _0861_/X vssd1 vssd1 vccd1 vccd1 _1600_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 hold382/X vssd1 vssd1 vccd1 vccd1 _0995_/C sky130_fd_sc_hd__clkbuf_2
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1510_ _1612_/CLK _1510_/D _1292_/Y vssd1 vssd1 vccd1 vccd1 _1510_/Q sky130_fd_sc_hd__dfrtp_1
X_1441_ _1634_/CLK hold19/X _1223_/Y vssd1 vssd1 vccd1 vccd1 _1441_/Q sky130_fd_sc_hd__dfrtp_1
X_1372_ _1413_/A vssd1 vssd1 vccd1 vccd1 _1372_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0957__D _1100_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0941_ _0967_/B _1180_/A vssd1 vssd1 vccd1 vccd1 _0946_/C sky130_fd_sc_hd__and2b_1
X_0872_ hold372/X hold16/X _0874_/S vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__mux2_1
XFILLER_0_50_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1355_ _1413_/A vssd1 vssd1 vccd1 vccd1 _1355_/Y sky130_fd_sc_hd__inv_2
X_1424_ _1505_/CLK _1424_/D _1206_/Y vssd1 vssd1 vccd1 vccd1 _1424_/Q sky130_fd_sc_hd__dfrtp_1
X_1286_ _1410_/A vssd1 vssd1 vccd1 vccd1 _1286_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_41_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1071_ _1192_/C _1137_/D _1071_/S vssd1 vssd1 vccd1 vccd1 _1497_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_1_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1140_ _1140_/A _1178_/S vssd1 vssd1 vccd1 vccd1 _1141_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_55_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0924_ _0887_/B _0915_/C _0917_/A vssd1 vssd1 vccd1 vccd1 _0925_/B sky130_fd_sc_hd__a21oi_1
X_0855_ _0855_/A _0855_/B vssd1 vssd1 vccd1 vccd1 _0855_/X sky130_fd_sc_hd__or2_1
X_0786_ _0847_/A _0786_/B vssd1 vssd1 vccd1 vccd1 _0786_/Y sky130_fd_sc_hd__nor2_1
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlygate4sd3_1
X_1407_ _1409_/A vssd1 vssd1 vccd1 vccd1 _1407_/Y sky130_fd_sc_hd__inv_2
X_1338_ _1339_/A vssd1 vssd1 vccd1 vccd1 _1338_/Y sky130_fd_sc_hd__inv_2
X_1269_ _1404_/A vssd1 vssd1 vccd1 vccd1 _1269_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_46_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0979__B _1007_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1123_ hold220/X hold224/X _1133_/S vssd1 vssd1 vccd1 vccd1 _1468_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_18_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1054_ hold286/X _1069_/S _1008_/X _1031_/C vssd1 vssd1 vccd1 vccd1 _1514_/D sky130_fd_sc_hd__a22o_1
X_0907_ _0902_/Y _0905_/X _0906_/X _0925_/A _0905_/A vssd1 vssd1 vccd1 vccd1 _0907_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_43_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0973__C_N _1191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0838_ _1606_/Q _0831_/B _0837_/X _0831_/A _0837_/A vssd1 vssd1 vccd1 vccd1 _0838_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__1091__S0 _1007_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0769_ _0806_/A _0803_/A _0817_/A _0813_/A vssd1 vssd1 vccd1 vccd1 _0773_/A sky130_fd_sc_hd__or4b_1
XANTENNA__0991__B1 _1103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1082__S0 _1100_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold329 _0934_/X vssd1 vssd1 vccd1 vccd1 _1568_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold307 _1570_/Q vssd1 vssd1 vccd1 vccd1 _0886_/A sky130_fd_sc_hd__buf_1
XFILLER_0_25_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold318 _0790_/X vssd1 vssd1 vccd1 vccd1 _1625_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1106_ _0995_/C hold333/X _1133_/S vssd1 vssd1 vccd1 vccd1 _1485_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_17_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1037_ hold72/X _1061_/A2 _1005_/B _1030_/X vssd1 vssd1 vccd1 vccd1 _1531_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_33_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0964__A0 _1100_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0992__B _1007_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold126 _1515_/Q vssd1 vssd1 vccd1 vccd1 hold126/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 _0975_/X vssd1 vssd1 vccd1 vccd1 _1017_/A sky130_fd_sc_hd__clkbuf_2
Xhold104 _1494_/Q vssd1 vssd1 vccd1 vccd1 hold104/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold159 _1058_/X vssd1 vssd1 vccd1 vccd1 _1510_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1586_ _1586_/CLK _1586_/D _1368_/Y vssd1 vssd1 vccd1 vccd1 _1586_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold137 _1557_/Q vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 _0991_/X vssd1 vssd1 vccd1 vccd1 _1552_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1371_ _1413_/A vssd1 vssd1 vccd1 vccd1 _1371_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_4_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1440_ _1624_/CLK _1440_/D _1222_/Y vssd1 vssd1 vccd1 vccd1 _1440_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1105__A0 _1191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1040__A2_N _1031_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1569_ _1583_/CLK _1569_/D _1351_/Y vssd1 vssd1 vccd1 vccd1 _1569_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0940_ input4/X _0939_/Y hold107/X _1101_/C vssd1 vssd1 vccd1 vccd1 _1179_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0871_ hold84/X hold208/X _0874_/S vssd1 vssd1 vccd1 vccd1 _0871_/X sky130_fd_sc_hd__mux2_1
X_1354_ _1413_/A vssd1 vssd1 vccd1 vccd1 _1354_/Y sky130_fd_sc_hd__inv_2
X_1423_ _1598_/CLK _1423_/D _1205_/Y vssd1 vssd1 vccd1 vccd1 _1423_/Q sky130_fd_sc_hd__dfrtp_2
X_1285_ _1410_/A vssd1 vssd1 vccd1 vccd1 _1285_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_41_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1020__A2 _1059_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1070_ _1007_/C _1187_/C _1071_/S vssd1 vssd1 vccd1 vccd1 _1498_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_55_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0923_ _0917_/Y _0922_/X _0923_/S vssd1 vssd1 vccd1 vccd1 _0923_/X sky130_fd_sc_hd__mux2_1
X_0854_ _0847_/A _0852_/X _0853_/X _0789_/A vssd1 vssd1 vccd1 vccd1 _0855_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_7_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0785_ _0786_/B _0784_/B _0783_/X vssd1 vssd1 vccd1 vccd1 _0785_/X sky130_fd_sc_hd__a21o_1
X_1337_ _1413_/A vssd1 vssd1 vccd1 vccd1 _1337_/Y sky130_fd_sc_hd__inv_2
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__dlygate4sd3_1
X_1268_ _1387_/A vssd1 vssd1 vccd1 vccd1 _1268_/Y sky130_fd_sc_hd__inv_2
X_1406_ _1409_/A vssd1 vssd1 vccd1 vccd1 _1406_/Y sky130_fd_sc_hd__inv_2
X_1199_ _0917_/A _1198_/Y _1595_/D vssd1 vssd1 vccd1 vccd1 _1566_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1122_ hold52/X _1469_/Q _1135_/S vssd1 vssd1 vccd1 vccd1 hold53/A sky130_fd_sc_hd__mux2_1
XANTENNA__0995__B _1100_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1053_ hold126/X _1061_/A2 _1005_/X _1031_/C vssd1 vssd1 vccd1 vccd1 _1053_/X sky130_fd_sc_hd__a22o_1
XANTENNA__1111__S _1133_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0906_ _0933_/B _0906_/B vssd1 vssd1 vccd1 vccd1 _0906_/X sky130_fd_sc_hd__and2_1
XFILLER_0_43_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0837_ _0837_/A _0837_/B vssd1 vssd1 vccd1 vccd1 _0837_/X sky130_fd_sc_hd__or2_1
XFILLER_0_22_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1091__S1 _1100_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0768_ _0850_/A _0768_/B vssd1 vssd1 vccd1 vccd1 _0786_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_11_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout105_A _1173_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1082__S1 _1100_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold308 _0929_/Y vssd1 vssd1 vccd1 vccd1 _1570_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold319 _1612_/Q vssd1 vssd1 vccd1 vccd1 _0837_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1105_ _1191_/B hold325/X _1133_/S vssd1 vssd1 vccd1 vccd1 _1486_/D sky130_fd_sc_hd__mux2_1
XANTENNA__1106__S _1133_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1036_ hold58/X _1061_/A2 _1002_/B _1030_/X vssd1 vssd1 vccd1 vccd1 hold59/A sky130_fd_sc_hd__a22o_1
XFILLER_0_31_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0992__C _1191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold127 _1053_/X vssd1 vssd1 vccd1 vccd1 _1515_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 _1538_/Q vssd1 vssd1 vccd1 vccd1 hold149/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 _0976_/X vssd1 vssd1 vccd1 vccd1 _1558_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 _0978_/X vssd1 vssd1 vccd1 vccd1 _1557_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold105 _1084_/X vssd1 vssd1 vccd1 vccd1 _1494_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1585_ _1586_/CLK _1585_/D _1367_/Y vssd1 vssd1 vccd1 vccd1 _1585_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1019_ _1019_/A _1027_/B vssd1 vssd1 vccd1 vccd1 _1019_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_8_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0873__A0 _1007_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1370_ _1413_/A vssd1 vssd1 vccd1 vccd1 _1370_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_45_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1568_ _1583_/CLK _1568_/D _1350_/Y vssd1 vssd1 vccd1 vccd1 _1568_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1499_ _1631_/CLK _1499_/D _1281_/Y vssd1 vssd1 vccd1 vccd1 _1499_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0870_ _1192_/D hold24/X _0874_/S vssd1 vssd1 vccd1 vccd1 _0870_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_50_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1422_ _1632_/CLK _1422_/D _1204_/Y vssd1 vssd1 vccd1 vccd1 _1636_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_0_2_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0998__B _1007_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1353_ _1413_/A vssd1 vssd1 vccd1 vccd1 _1353_/Y sky130_fd_sc_hd__inv_2
X_1284_ _1387_/A vssd1 vssd1 vccd1 vccd1 _1284_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1114__S _1133_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1014__B1 _0970_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0999_ hold81/X _0999_/B vssd1 vssd1 vccd1 vccd1 _0999_/X sky130_fd_sc_hd__and2_1
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0922_ _0917_/B _0906_/X _0925_/A vssd1 vssd1 vccd1 vccd1 _0922_/X sky130_fd_sc_hd__a21o_1
X_0853_ hold48/X _1598_/Q hold62/X _1602_/Q _0851_/S _0850_/A vssd1 vssd1 vccd1 vccd1
+ _0853_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_46_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1405_ _1405_/A vssd1 vssd1 vccd1 vccd1 _1405_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_23_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0784_ _0786_/B _0784_/B vssd1 vssd1 vccd1 vccd1 _0784_/X sky130_fd_sc_hd__and2_1
XANTENNA__1109__S _1133_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput1 i_start_rx vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1198_ hold30/X input1/X vssd1 vssd1 vccd1 vccd1 _1198_/Y sky130_fd_sc_hd__nand2b_1
X_1336_ _1417_/A vssd1 vssd1 vccd1 vccd1 _1336_/Y sky130_fd_sc_hd__inv_2
X_1267_ _1339_/A vssd1 vssd1 vccd1 vccd1 _1267_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_46_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1052_ hold265/X _1071_/S _1002_/X _1031_/C vssd1 vssd1 vccd1 vccd1 _1516_/D sky130_fd_sc_hd__a22o_1
XANTENNA__0995__C _0995_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1121_ hold76/X _1470_/Q _1133_/S vssd1 vssd1 vccd1 vccd1 hold77/A sky130_fd_sc_hd__mux2_1
XANTENNA__0986__A1_N _0971_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0905_ _0905_/A _0905_/B vssd1 vssd1 vccd1 vccd1 _0905_/X sky130_fd_sc_hd__or2_1
XFILLER_0_43_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0836_ _0836_/A _0836_/B _0836_/C vssd1 vssd1 vccd1 vccd1 _1613_/D sky130_fd_sc_hd__and3_1
XFILLER_0_28_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0767_ _0789_/A _0851_/S vssd1 vssd1 vccd1 vccd1 _0767_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_11_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0991__A2 _1069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1319_ _1404_/A vssd1 vssd1 vccd1 vccd1 _1319_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_2_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold309 _1614_/Q vssd1 vssd1 vccd1 vccd1 _0833_/A sky130_fd_sc_hd__buf_1
XFILLER_0_33_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1122__S _1135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1104_ _0989_/C hold269/X _1135_/S vssd1 vssd1 vccd1 vccd1 _1487_/D sky130_fd_sc_hd__mux2_1
X_1035_ hold98/X _1071_/S _0999_/B _1030_/X vssd1 vssd1 vccd1 vccd1 _1035_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_16_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0819_ _0803_/A _0820_/B _0818_/Y vssd1 vssd1 vccd1 vccd1 _0819_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_19_clk_A clkbuf_1_1__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1584_ _1635_/CLK _1584_/D _1366_/Y vssd1 vssd1 vccd1 vccd1 _1584_/Q sky130_fd_sc_hd__dfrtp_1
Xhold139 _1635_/Q vssd1 vssd1 vccd1 vccd1 hold139/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold106 _1421_/Q vssd1 vssd1 vccd1 vccd1 _1101_/B sky130_fd_sc_hd__buf_1
Xhold128 hold380/X vssd1 vssd1 vccd1 vccd1 _1192_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_0_0_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold117 hold379/X vssd1 vssd1 vccd1 vccd1 _1192_/C sky130_fd_sc_hd__clkbuf_2
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1117__S _1135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1018_ hold154/X _1059_/A2 _1103_/B _1017_/Y vssd1 vssd1 vccd1 vccd1 _1018_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_44_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1050__B2 _1031_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1636_ _1636_/A vssd1 vssd1 vccd1 vccd1 _1636_/X sky130_fd_sc_hd__clkbuf_2
X_1567_ _1582_/CLK _1567_/D _1349_/Y vssd1 vssd1 vccd1 vccd1 _1567_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1041__B2 _1059_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1498_ _1631_/CLK _1498_/D _1280_/Y vssd1 vssd1 vccd1 vccd1 _1498_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1032__B2 _1030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1421_ _1625_/CLK _1421_/D _1203_/Y vssd1 vssd1 vccd1 vccd1 _1421_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_2_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1352_ _1363_/A vssd1 vssd1 vccd1 vccd1 _1352_/Y sky130_fd_sc_hd__inv_2
X_1283_ _1410_/A vssd1 vssd1 vccd1 vccd1 _1283_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1130__S _1135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout128_A _1416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0998_ _1100_/A _1007_/B _1192_/D vssd1 vssd1 vccd1 vccd1 _0999_/B sky130_fd_sc_hd__and3b_1
X_1619_ _1627_/CLK _1619_/D _1401_/Y vssd1 vssd1 vccd1 vccd1 _1619_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0921_ _0921_/A vssd1 vssd1 vccd1 vccd1 _1574_/D sky130_fd_sc_hd__inv_2
XFILLER_0_55_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0783_ _0826_/B _0782_/B _0831_/A vssd1 vssd1 vccd1 vccd1 _0783_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_11_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0852_ _0852_/A _0852_/B vssd1 vssd1 vccd1 vccd1 _0852_/X sky130_fd_sc_hd__or2_1
X_1404_ _1404_/A vssd1 vssd1 vccd1 vccd1 _1404_/Y sky130_fd_sc_hd__inv_2
X_1335_ _1384_/A vssd1 vssd1 vccd1 vccd1 _1335_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_39_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput2 i_uart_rx vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1125__S _1133_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1266_ _1415_/A vssd1 vssd1 vccd1 vccd1 _1266_/Y sky130_fd_sc_hd__inv_2
X_1197_ hold277/X _1183_/Y _1196_/X _1183_/B _1180_/A vssd1 vssd1 vccd1 vccd1 _1418_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_46_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0994__B1 _1103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1094__S0 _1100_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1085__S0 _1100_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1120_ hold147/X hold188/X _1133_/S vssd1 vssd1 vccd1 vccd1 _1120_/X sky130_fd_sc_hd__mux2_1
X_1051_ hold34/X _1069_/S _0999_/X _1031_/C vssd1 vssd1 vccd1 vccd1 _1517_/D sky130_fd_sc_hd__a22o_1
X_0904_ _1566_/Q _0894_/Y _0903_/X _0925_/A _0893_/A vssd1 vssd1 vccd1 vccd1 _0904_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_28_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0835_ _0835_/A _0835_/B vssd1 vssd1 vccd1 vccd1 _0836_/C sky130_fd_sc_hd__or2_1
XANTENNA__1076__S0 _1100_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0766_ _0789_/A _1624_/Q vssd1 vssd1 vccd1 vccd1 _0766_/X sky130_fd_sc_hd__and2_1
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1318_ _1339_/A vssd1 vssd1 vccd1 vccd1 _1318_/Y sky130_fd_sc_hd__inv_2
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1249_ _1404_/A vssd1 vssd1 vccd1 vccd1 _1249_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_19_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1034_ hold253/X _1061_/A2 _0996_/B _1030_/X vssd1 vssd1 vccd1 vccd1 _1534_/D sky130_fd_sc_hd__a22o_1
X_1103_ _1178_/S _1103_/B vssd1 vssd1 vccd1 vccd1 _1129_/S sky130_fd_sc_hd__nand2_4
X_0749_ _0753_/D hold55/X vssd1 vssd1 vccd1 vccd1 hold56/A sky130_fd_sc_hd__nor2_1
X_0818_ _0803_/A _0820_/B _0836_/A vssd1 vssd1 vccd1 vccd1 _0818_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout110_A _0970_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1583_ _1583_/CLK _1583_/D _1365_/Y vssd1 vssd1 vccd1 vccd1 _1583_/Q sky130_fd_sc_hd__dfrtp_1
Xhold129 _0977_/X vssd1 vssd1 vccd1 vccd1 _1019_/A sky130_fd_sc_hd__buf_1
XFILLER_0_21_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold118 _1027_/A vssd1 vssd1 vccd1 vccd1 hold118/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold107 _0938_/Y vssd1 vssd1 vccd1 vccd1 hold107/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1108__A0 hold84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1133__S _1133_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1017_ _1017_/A _1027_/B vssd1 vssd1 vccd1 vccd1 _1017_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__1001__A_N _1100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1050__A2 _1059_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1128__S _1129_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1566_ _1589_/CLK _1566_/D _1348_/Y vssd1 vssd1 vccd1 vccd1 _1566_/Q sky130_fd_sc_hd__dfrtp_1
X_1635_ _1635_/CLK _1635_/D _1417_/Y vssd1 vssd1 vccd1 vccd1 _1635_/Q sky130_fd_sc_hd__dfrtp_1
X_1497_ _1631_/CLK _1497_/D _1279_/Y vssd1 vssd1 vccd1 vccd1 _1497_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_18_clk_A clkbuf_1_1__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1032__A2 _1069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1351_ _1363_/A vssd1 vssd1 vccd1 vccd1 _1351_/Y sky130_fd_sc_hd__inv_2
X_1420_ _1602_/CLK _1420_/D _1202_/Y vssd1 vssd1 vccd1 vccd1 _1420_/Q sky130_fd_sc_hd__dfrtp_1
X_1282_ _1410_/A vssd1 vssd1 vccd1 vccd1 _1282_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1191__B _1191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0997_ hold52/X _1061_/A2 _1103_/B _0996_/X vssd1 vssd1 vccd1 vccd1 _0997_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_41_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1618_ _1625_/CLK _1618_/D _1400_/Y vssd1 vssd1 vccd1 vccd1 _1618_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1549_ _1605_/CLK _1549_/D _1331_/Y vssd1 vssd1 vccd1 vccd1 _1549_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold290 _0914_/X vssd1 vssd1 vccd1 vccd1 _1576_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0920_ _0919_/Y _0919_/A _0920_/S vssd1 vssd1 vccd1 vccd1 _0921_/A sky130_fd_sc_hd__mux2_1
X_0782_ _1606_/Q _0782_/B vssd1 vssd1 vccd1 vccd1 _0782_/X sky130_fd_sc_hd__and2_1
XFILLER_0_11_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0851_ _1603_/Q hold12/X _0851_/S vssd1 vssd1 vccd1 vccd1 _0852_/B sky130_fd_sc_hd__mux2_1
X_1265_ _1363_/A vssd1 vssd1 vccd1 vccd1 _1265_/Y sky130_fd_sc_hd__inv_2
X_1403_ _1409_/A vssd1 vssd1 vccd1 vccd1 _1403_/Y sky130_fd_sc_hd__inv_2
X_1334_ _1339_/A vssd1 vssd1 vccd1 vccd1 _1334_/Y sky130_fd_sc_hd__inv_2
Xinput3 rst vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_1
XFILLER_0_52_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1196_ _1187_/X _1188_/X _1184_/B vssd1 vssd1 vccd1 vccd1 _1196_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_52_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1094__S1 _1100_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1085__S1 _1100_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1050_ hold46/X _1059_/A2 _0996_/X _1031_/C vssd1 vssd1 vccd1 vccd1 _1518_/D sky130_fd_sc_hd__a22o_1
X_0903_ _1579_/Q _0905_/B _0893_/A vssd1 vssd1 vccd1 vccd1 _0903_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_43_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0834_ _0833_/A _0783_/X _0831_/X _0833_/Y vssd1 vssd1 vccd1 vccd1 _0834_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0976__B2 _1069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0765_ _0744_/X hold40/X _0765_/S vssd1 vssd1 vccd1 vccd1 _0765_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1076__S1 _1100_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1317_ _1415_/A vssd1 vssd1 vccd1 vccd1 _1317_/Y sky130_fd_sc_hd__inv_2
X_1248_ _1385_/A vssd1 vssd1 vccd1 vccd1 _1248_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_2_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1179_ _1179_/A _1179_/B _1179_/C vssd1 vssd1 vccd1 vccd1 _1183_/B sky130_fd_sc_hd__or3_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1102_ _0775_/A _1073_/Y _1179_/B vssd1 vssd1 vccd1 vccd1 _1102_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1033_ hold236/X _1069_/S _0993_/B _1030_/X vssd1 vssd1 vccd1 vccd1 _1535_/D sky130_fd_sc_hd__a22o_1
X_0817_ _0817_/A _1617_/Q _1606_/Q _0817_/D vssd1 vssd1 vccd1 vccd1 _0820_/B sky130_fd_sc_hd__and4_1
XFILLER_0_16_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0748_ _0753_/A _0880_/A vssd1 vssd1 vccd1 vccd1 hold55/A sky130_fd_sc_hd__or2_1
XFILLER_0_39_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1053__B1 _1005_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold108 _1096_/S vssd1 vssd1 vccd1 vccd1 _1099_/S sky130_fd_sc_hd__buf_2
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1582_ _1582_/CLK _1582_/D _1364_/Y vssd1 vssd1 vccd1 vccd1 _1582_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold119 _0986_/X vssd1 vssd1 vccd1 vccd1 _1553_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1016_ hold110/X _1061_/A2 _0970_/X _1015_/Y vssd1 vssd1 vccd1 vccd1 _1016_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_8_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_20_clk clkbuf_1_1__f_clk/X vssd1 vssd1 vccd1 vccd1 _1601_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_45_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_11_clk clkbuf_1_1__f_clk/X vssd1 vssd1 vccd1 vccd1 _1544_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__1026__B1 _1103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1634_ _1634_/CLK hold57/X _1416_/Y vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__1144__S _1168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1565_ _1624_/CLK input2/X _1347_/Y vssd1 vssd1 vccd1 vccd1 _1565_/Q sky130_fd_sc_hd__dfstp_1
X_1496_ _1547_/CLK _1496_/D _1278_/Y vssd1 vssd1 vccd1 vccd1 _1496_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0984__A1_N _0971_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1350_ _1363_/A vssd1 vssd1 vccd1 vccd1 _1350_/Y sky130_fd_sc_hd__inv_2
X_1281_ _1410_/A vssd1 vssd1 vccd1 vccd1 _1281_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_0_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _1556_/CLK sky130_fd_sc_hd__clkbuf_16
X_0996_ hold81/X _0996_/B vssd1 vssd1 vccd1 vccd1 _0996_/X sky130_fd_sc_hd__and2_1
XFILLER_0_41_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1617_ _1627_/CLK _1617_/D _1399_/Y vssd1 vssd1 vccd1 vccd1 _1617_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1479_ _1544_/CLK _1479_/D _1261_/Y vssd1 vssd1 vccd1 vccd1 _1479_/Q sky130_fd_sc_hd__dfrtp_1
X_1548_ _1548_/CLK hold85/X _1330_/Y vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold280 _1182_/X vssd1 vssd1 vccd1 vccd1 _1421_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 _1625_/Q vssd1 vssd1 vccd1 vccd1 _0789_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0850_ _0850_/A _1625_/Q vssd1 vssd1 vccd1 vccd1 _0850_/X sky130_fd_sc_hd__or2_1
X_0781_ _0781_/A _0781_/B _0781_/C _0781_/D vssd1 vssd1 vccd1 vccd1 _0782_/B sky130_fd_sc_hd__or4_1
X_1402_ _1402_/A vssd1 vssd1 vccd1 vccd1 _1402_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_23_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_17_clk_A clkbuf_1_1__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1333_ _1415_/A vssd1 vssd1 vccd1 vccd1 _1333_/Y sky130_fd_sc_hd__inv_2
X_1264_ _1384_/A vssd1 vssd1 vccd1 vccd1 _1264_/Y sky130_fd_sc_hd__inv_2
Xinput4 wb_ack_i vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_1
X_1195_ _0967_/B _1183_/B _1183_/Y _1194_/X vssd1 vssd1 vccd1 vccd1 _1419_/D sky130_fd_sc_hd__a22o_1
X_0979_ _1100_/A _1007_/B hold84/X vssd1 vssd1 vccd1 vccd1 _1021_/A sky130_fd_sc_hd__or3b_2
XFILLER_0_14_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0994__A2 _1069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0902_ _0905_/A _0905_/B vssd1 vssd1 vccd1 vccd1 _0902_/Y sky130_fd_sc_hd__nand2_1
X_0833_ _0833_/A _0836_/B vssd1 vssd1 vccd1 vccd1 _0833_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_22_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0764_ _0764_/A _0764_/B _0764_/C _0764_/D vssd1 vssd1 vccd1 vccd1 _0764_/X sky130_fd_sc_hd__or4_1
XFILLER_0_11_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1316_ _1405_/A vssd1 vssd1 vccd1 vccd1 _1316_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_2_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1152__S _1168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1247_ _1415_/A vssd1 vssd1 vccd1 vccd1 _1247_/Y sky130_fd_sc_hd__inv_2
X_1178_ _1031_/C _1141_/C _1178_/S vssd1 vssd1 vccd1 vccd1 _1180_/B sky130_fd_sc_hd__mux2_1
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1101_ _0775_/A _1101_/B _1101_/C _1101_/D vssd1 vssd1 vccd1 vccd1 _1179_/B sky130_fd_sc_hd__and4b_1
X_1032_ hold234/X _1069_/S hold144/X _1030_/X vssd1 vssd1 vccd1 vccd1 _1536_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_33_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0747_ _0764_/A _0884_/S vssd1 vssd1 vccd1 vccd1 _0880_/A sky130_fd_sc_hd__nand2_1
XANTENNA__1147__S _1173_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0816_ _0822_/A _1606_/Q _0817_/D vssd1 vssd1 vccd1 vccd1 _0816_/X sky130_fd_sc_hd__and3_1
XFILLER_0_3_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1062__B2 _1031_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1581_ _1582_/CLK _1581_/D _1363_/Y vssd1 vssd1 vccd1 vccd1 _1581_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1053__B2 _1031_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold109 _1081_/X vssd1 vssd1 vccd1 vccd1 _1495_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1015_ _1015_/A _1027_/B vssd1 vssd1 vccd1 vccd1 _1015_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_56_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1044__B2 _1071_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0979__C_N hold84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1035__B2 _1030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1633_ _1635_/CLK hold31/X _1415_/Y vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__dfrtp_1
X_1564_ _1605_/CLK _1564_/D _1346_/Y vssd1 vssd1 vccd1 vccd1 _1564_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1495_ _1600_/CLK _1495_/D _1277_/Y vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__dfrtp_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1160__S _1168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1070__S _1071_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1280_ _1413_/A vssd1 vssd1 vccd1 vccd1 _1280_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_25_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0995_ _0981_/A _1100_/C _0995_/C vssd1 vssd1 vccd1 vccd1 _0996_/B sky130_fd_sc_hd__and3b_1
XFILLER_0_26_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1155__S _1168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1616_ _1627_/CLK _1616_/D _1398_/Y vssd1 vssd1 vccd1 vccd1 _1616_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1547_ _1547_/CLK _1547_/D _1329_/Y vssd1 vssd1 vccd1 vccd1 _1547_/Q sky130_fd_sc_hd__dfrtp_1
X_1478_ _1544_/CLK hold45/X _1260_/Y vssd1 vssd1 vccd1 vccd1 _1478_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_49_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0997__B1 _1103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1097__S0 _1007_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold281 _1575_/Q vssd1 vssd1 vccd1 vccd1 _0912_/A sky130_fd_sc_hd__buf_1
Xhold270 _1611_/Q vssd1 vssd1 vccd1 vccd1 _0795_/A sky130_fd_sc_hd__buf_1
Xhold292 _0766_/X vssd1 vssd1 vccd1 vccd1 _0768_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1065__S _1071_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0780_ _0780_/A _0807_/A _0806_/A _0813_/A vssd1 vssd1 vccd1 vccd1 _0781_/D sky130_fd_sc_hd__or4b_1
XANTENNA__1088__S0 _1100_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1401_ _1409_/A vssd1 vssd1 vccd1 vccd1 _1401_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_11_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput5 wb_dat_i[0] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_1
X_1332_ _1405_/A vssd1 vssd1 vccd1 vccd1 _1332_/Y sky130_fd_sc_hd__inv_2
X_1263_ _1405_/A vssd1 vssd1 vccd1 vccd1 _1263_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_39_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1194_ _0995_/C _1007_/C _1073_/B _1193_/X _1189_/X vssd1 vssd1 vccd1 vccd1 _1194_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout126_A _1416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0978_ _0971_/Y _0977_/X hold38/X _1069_/S vssd1 vssd1 vccd1 vccd1 _0978_/X sky130_fd_sc_hd__a2bb2o_1
XANTENNA__1079__S0 _1100_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0901_ _0933_/B _0895_/Y _0900_/X _0925_/A _0896_/A vssd1 vssd1 vccd1 vccd1 _0901_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_51_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0832_ _0835_/A _0835_/B vssd1 vssd1 vccd1 vccd1 _0836_/B sky130_fd_sc_hd__nand2_1
X_0763_ _0764_/A _0764_/B hold30/X _0758_/Y _0762_/X vssd1 vssd1 vccd1 vccd1 _1629_/D
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_11_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1315_ _1387_/A vssd1 vssd1 vccd1 vccd1 _1315_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_37_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1177_ hold272/X _1176_/X _1135_/S vssd1 vssd1 vccd1 vccd1 _1177_/X sky130_fd_sc_hd__a21bo_1
X_1246_ _1384_/A vssd1 vssd1 vccd1 vccd1 _1246_/Y sky130_fd_sc_hd__inv_2
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_16_clk_A clkbuf_1_1__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1031_ hold86/X _1100_/B _1031_/C vssd1 vssd1 vccd1 vccd1 _1031_/Y sky130_fd_sc_hd__nand3b_4
X_1100_ _1100_/A _1100_/B _1100_/C hold86/X vssd1 vssd1 vccd1 vccd1 _1101_/D sky130_fd_sc_hd__or4b_1
XFILLER_0_56_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1001__B _1100_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0746_ hold30/X _0882_/B _0745_/X _0742_/X vssd1 vssd1 vccd1 vccd1 _1635_/D sky130_fd_sc_hd__a31o_1
X_0815_ _1606_/Q _0817_/D vssd1 vssd1 vccd1 vccd1 _0825_/B sky130_fd_sc_hd__nand2_1
Xinput30 wb_dat_i[3] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__buf_1
XANTENNA__1163__S _1168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1229_ _1397_/A vssd1 vssd1 vccd1 vccd1 _1229_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_53_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1580_ _1580_/CLK _1580_/D _1362_/Y vssd1 vssd1 vccd1 vccd1 _1580_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1014_ hold259/X _1061_/A2 _0970_/X _1013_/Y vssd1 vssd1 vccd1 vccd1 _1544_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_44_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1158__S _1173_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0729_ _0893_/A _0892_/A _0892_/B _0905_/A vssd1 vssd1 vccd1 vccd1 _0740_/A sky130_fd_sc_hd__or4b_1
XFILLER_0_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1035__A2 _1071_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1026__A2 _1071_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1632_ _1632_/CLK hold25/X _1414_/Y vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__dfrtp_1
X_1494_ _1601_/CLK _1494_/D _1276_/Y vssd1 vssd1 vccd1 vccd1 _1494_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1563_ _1600_/CLK _1563_/D _1345_/Y vssd1 vssd1 vccd1 vccd1 _1563_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0994_ hold76/X _1069_/S _1103_/B hold82/X vssd1 vssd1 vccd1 vccd1 hold83/A sky130_fd_sc_hd__a22o_1
XFILLER_0_14_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1615_ _1615_/CLK _1615_/D _1397_/Y vssd1 vssd1 vccd1 vccd1 _1615_/Q sky130_fd_sc_hd__dfrtp_1
X_1477_ _1558_/CLK hold67/X _1259_/Y vssd1 vssd1 vccd1 vccd1 _1477_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1546_ _1556_/CLK hold91/X _1328_/Y vssd1 vssd1 vccd1 vccd1 hold90/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1171__S _1171_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold260 _1128_/X vssd1 vssd1 vccd1 vccd1 _1463_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 _0840_/X vssd1 vssd1 vccd1 vccd1 _1611_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1097__S1 _1100_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold282 _0916_/X vssd1 vssd1 vccd1 vccd1 _1575_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 _0788_/X vssd1 vssd1 vccd1 vccd1 _1626_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1088__S1 _1100_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1400_ _1409_/A vssd1 vssd1 vccd1 vccd1 _1400_/Y sky130_fd_sc_hd__inv_2
X_1331_ _1387_/A vssd1 vssd1 vccd1 vccd1 _1331_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput6 wb_dat_i[10] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__buf_1
XANTENNA__1004__B _1100_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1193_ _1191_/A _1191_/B _1192_/X _1191_/Y vssd1 vssd1 vccd1 vccd1 _1193_/X sky130_fd_sc_hd__a31o_1
X_1262_ _1387_/A vssd1 vssd1 vccd1 vccd1 _1262_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_52_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0977_ _1100_/A _1007_/B _1192_/D vssd1 vssd1 vccd1 vccd1 _0977_/X sky130_fd_sc_hd__or3b_2
XANTENNA__1166__S _1168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1079__S1 _1100_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout119_A _1416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1529_ _1548_/CLK _1529_/D _1311_/Y vssd1 vssd1 vccd1 vccd1 _1529_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0900_ _0905_/B _0896_/D _0896_/A vssd1 vssd1 vccd1 vccd1 _0900_/X sky130_fd_sc_hd__a21o_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0831_ _0831_/A _0831_/B _1613_/Q vssd1 vssd1 vccd1 vccd1 _0831_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_36_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0762_ _0754_/A _0884_/S _0753_/D _0758_/B hold210/X vssd1 vssd1 vccd1 vccd1 _0762_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1314_ _1404_/A vssd1 vssd1 vccd1 vccd1 _1314_/Y sky130_fd_sc_hd__inv_2
X_1245_ _1363_/A vssd1 vssd1 vccd1 vccd1 _1245_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1015__A _1015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1176_ _1140_/A _1178_/S _1141_/C _1179_/C _1175_/X vssd1 vssd1 vccd1 vccd1 _1176_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_34_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0982__A1_N _0971_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1065__A0 _1191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1030_ hold86/X _1100_/B _1031_/C vssd1 vssd1 vccd1 vccd1 _1030_/X sky130_fd_sc_hd__and3b_4
XANTENNA__1001__C hold84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput20 wb_dat_i[23] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__buf_1
X_0814_ _0782_/X _0805_/Y _0813_/X _0831_/A _0813_/A vssd1 vssd1 vccd1 vccd1 _0814_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_3_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput31 wb_dat_i[4] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__buf_1
X_0745_ _0764_/D _0758_/B vssd1 vssd1 vccd1 vccd1 _0745_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1228_ _1385_/A vssd1 vssd1 vccd1 vccd1 _1228_/Y sky130_fd_sc_hd__inv_2
X_1159_ hold202/X _1438_/Q _1173_/S vssd1 vssd1 vccd1 vccd1 _1159_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_30_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0989__A_N _1100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_23_clk clkbuf_1_1__f_clk/X vssd1 vssd1 vccd1 vccd1 _1489_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1013_ _1013_/A _1027_/B vssd1 vssd1 vccd1 vccd1 _1013_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_56_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_14_clk clkbuf_1_1__f_clk/X vssd1 vssd1 vccd1 vccd1 _1623_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_8_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0728_ _0741_/C vssd1 vssd1 vccd1 vccd1 _0866_/A sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_15_clk_A clkbuf_1_1__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1631_ _1631_/CLK _1631_/D _1413_/Y vssd1 vssd1 vccd1 vccd1 _1631_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_3_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _1631_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1562_ _1562_/CLK _1562_/D _1344_/Y vssd1 vssd1 vccd1 vccd1 hold80/A sky130_fd_sc_hd__dfrtp_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1493_ _1600_/CLK _1493_/D _1275_/Y vssd1 vssd1 vccd1 vccd1 _1493_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1007__B _1007_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1169__S _1171_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0993_ hold81/X _0993_/B vssd1 vssd1 vccd1 vccd1 hold82/A sky130_fd_sc_hd__and2_1
XFILLER_0_41_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1614_ _1615_/CLK _1614_/D _1396_/Y vssd1 vssd1 vccd1 vccd1 _1614_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1476_ _1558_/CLK hold39/X _1258_/Y vssd1 vssd1 vccd1 vccd1 _1476_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1545_ _1601_/CLK _1545_/D _1327_/Y vssd1 vssd1 vccd1 vccd1 _1545_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold261 _1566_/Q vssd1 vssd1 vccd1 vccd1 _0933_/B sky130_fd_sc_hd__clkbuf_4
Xhold294 _1583_/Q vssd1 vssd1 vccd1 vccd1 _0884_/S sky130_fd_sc_hd__buf_2
Xhold272 _1423_/Q vssd1 vssd1 vccd1 vccd1 hold272/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 _1418_/Q vssd1 vssd1 vccd1 vccd1 _1180_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold250 _1454_/Q vssd1 vssd1 vccd1 vccd1 hold250/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1261_ _1405_/A vssd1 vssd1 vccd1 vccd1 _1261_/Y sky130_fd_sc_hd__inv_2
X_1330_ _1404_/A vssd1 vssd1 vccd1 vccd1 _1330_/Y sky130_fd_sc_hd__inv_2
X_1192_ _1590_/Q _1192_/B _1192_/C _1192_/D vssd1 vssd1 vccd1 vccd1 _1192_/X sky130_fd_sc_hd__and4b_1
Xinput7 wb_dat_i[11] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_1
XFILLER_0_54_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0976_ _0971_/Y _0975_/X hold66/X _1069_/S vssd1 vssd1 vccd1 vccd1 _0976_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_6_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1528_ _1623_/CLK _1528_/D _1310_/Y vssd1 vssd1 vccd1 vccd1 _1528_/Q sky130_fd_sc_hd__dfrtp_1
X_1459_ _1605_/CLK _1459_/D _1241_/Y vssd1 vssd1 vccd1 vccd1 _1459_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0830_ _0830_/A vssd1 vssd1 vccd1 vccd1 _1615_/D sky130_fd_sc_hd__inv_2
XFILLER_0_22_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0761_ _0764_/A _0884_/S hold30/X _0758_/Y _0760_/X vssd1 vssd1 vccd1 vccd1 _0761_/X
+ sky130_fd_sc_hd__a41o_1
X_1244_ _1405_/A vssd1 vssd1 vccd1 vccd1 _1244_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1313_ _1404_/A vssd1 vssd1 vccd1 vccd1 _1313_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1015__B _1027_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1175_ _0720_/Y _0939_/Y _0946_/C _1420_/Q vssd1 vssd1 vccd1 vccd1 _1175_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_42_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0959_ _1100_/B _1100_/C hold86/X vssd1 vssd1 vccd1 vccd1 _0960_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_33_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0813_ _0813_/A _0813_/B vssd1 vssd1 vccd1 vccd1 _0813_/X sky130_fd_sc_hd__or2_1
Xinput21 wb_dat_i[24] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput10 wb_dat_i[14] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__buf_1
Xinput32 wb_dat_i[5] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1056__B2 _1031_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0744_ _0726_/A _0764_/C hold30/X vssd1 vssd1 vccd1 vccd1 _0744_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_42_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1158_ hold100/X _1439_/Q _1173_/S vssd1 vssd1 vccd1 vccd1 _1158_/X sky130_fd_sc_hd__mux2_1
X_1227_ _1385_/A vssd1 vssd1 vccd1 vccd1 _1227_/Y sky130_fd_sc_hd__inv_2
X_1089_ _1098_/A _1089_/B vssd1 vssd1 vccd1 vccd1 _1089_/X sky130_fd_sc_hd__and2_1
XANTENNA__1047__B2 _1059_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1038__B2 _1030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1012_ hold171/X _1059_/A2 _1103_/B _1011_/X vssd1 vssd1 vccd1 vccd1 _1545_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0727_ hold54/X _0726_/A _0882_/A vssd1 vssd1 vccd1 vccd1 _0741_/C sky130_fd_sc_hd__o21a_1
XFILLER_0_8_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1630_ _1631_/CLK _1630_/D _1412_/Y vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1007__C _1007_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1492_ _1547_/CLK _1492_/D _1274_/Y vssd1 vssd1 vccd1 vccd1 _1492_/Q sky130_fd_sc_hd__dfrtp_1
X_1561_ _1562_/CLK _1561_/D _1343_/Y vssd1 vssd1 vccd1 vccd1 hold94/A sky130_fd_sc_hd__dfrtp_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1023__B _1027_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1110__A0 _1007_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_14_clk_A clkbuf_1_1__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0992_ _1100_/A _1007_/B _1191_/B vssd1 vssd1 vccd1 vccd1 _0993_/B sky130_fd_sc_hd__and3b_1
X_1544_ _1544_/CLK _1544_/D _1326_/Y vssd1 vssd1 vccd1 vccd1 _1544_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1613_ _1615_/CLK _1613_/D _1395_/Y vssd1 vssd1 vccd1 vccd1 _1613_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1475_ _1556_/CLK hold23/X _1257_/Y vssd1 vssd1 vccd1 vccd1 _1475_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1007__A_N _1564_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold295 _0761_/X vssd1 vssd1 vccd1 vccd1 _1630_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 _0878_/X vssd1 vssd1 vccd1 vccd1 hold262/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 _1610_/Q vssd1 vssd1 vccd1 vccd1 _0795_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold240 _1150_/X vssd1 vssd1 vccd1 vccd1 _1447_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 _1177_/X vssd1 vssd1 vccd1 vccd1 _1423_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 _1143_/X vssd1 vssd1 vccd1 vccd1 _1454_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1260_ _1405_/A vssd1 vssd1 vccd1 vccd1 _1260_/Y sky130_fd_sc_hd__inv_2
X_1191_ _1191_/A _1191_/B _1191_/C vssd1 vssd1 vccd1 vccd1 _1191_/Y sky130_fd_sc_hd__nor3_1
Xinput8 wb_dat_i[12] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_1
XFILLER_0_52_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0975_ _1100_/A _1007_/B _0995_/C vssd1 vssd1 vccd1 vccd1 _0975_/X sky130_fd_sc_hd__or3b_2
X_1527_ _1547_/CLK _1527_/D _1309_/Y vssd1 vssd1 vccd1 vccd1 hold70/A sky130_fd_sc_hd__dfrtp_1
X_1389_ _1402_/A vssd1 vssd1 vccd1 vccd1 _1389_/Y sky130_fd_sc_hd__inv_2
X_1458_ _1605_/CLK _1458_/D _1240_/Y vssd1 vssd1 vccd1 vccd1 _1458_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0760_ _0764_/C _0753_/D _0880_/A hold16/X vssd1 vssd1 vccd1 vccd1 _0760_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_36_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1243_ _1397_/A vssd1 vssd1 vccd1 vccd1 _1243_/Y sky130_fd_sc_hd__inv_2
X_1312_ _1417_/A vssd1 vssd1 vccd1 vccd1 _1312_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_2_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1174_ _1140_/A _1178_/S _1141_/A _1141_/B vssd1 vssd1 vccd1 vccd1 _1179_/C sky130_fd_sc_hd__a211oi_1
XANTENNA__1031__B _1100_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0889_ _1574_/Q _0923_/S _0889_/C _1571_/Q vssd1 vssd1 vccd1 vccd1 _0915_/D sky130_fd_sc_hd__and4_1
XFILLER_0_42_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0958_ _1101_/C _1185_/B _1178_/S vssd1 vssd1 vccd1 vccd1 _0960_/C sky130_fd_sc_hd__or3b_1
XFILLER_0_10_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1056__A2 _1059_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput22 wb_dat_i[25] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__buf_1
Xinput11 wb_dat_i[15] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__buf_1
Xinput33 wb_dat_i[6] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__clkbuf_2
X_0743_ hold54/X _0764_/A vssd1 vssd1 vccd1 vccd1 _0758_/B sky130_fd_sc_hd__xnor2_1
X_0812_ _0812_/A _0812_/B vssd1 vssd1 vccd1 vccd1 _1621_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_24_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_9_clk/A sky130_fd_sc_hd__clkbuf_16
X_1226_ _1397_/A vssd1 vssd1 vccd1 vccd1 _1226_/Y sky130_fd_sc_hd__inv_2
X_1157_ hold216/X _1440_/Q _1168_/S vssd1 vssd1 vccd1 vccd1 _1157_/X sky130_fd_sc_hd__mux2_1
X_1088_ input30/X input7/X input15/X input24/X _1100_/C _1100_/B vssd1 vssd1 vccd1
+ vccd1 _1089_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_30_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1038__A2 _1071_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1011_ hold81/X _1011_/B vssd1 vssd1 vccd1 vccd1 _1011_/X sky130_fd_sc_hd__and2_1
XFILLER_0_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0726_ _0726_/A _0764_/C vssd1 vssd1 vccd1 vccd1 _0741_/B sky130_fd_sc_hd__nor2_1
X_1209_ _1339_/A vssd1 vssd1 vccd1 vccd1 _1209_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_50_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1560_ _1623_/CLK _1560_/D _1342_/Y vssd1 vssd1 vccd1 vccd1 _1560_/Q sky130_fd_sc_hd__dfrtp_1
X_1491_ _1598_/CLK _1491_/D _1273_/Y vssd1 vssd1 vccd1 vccd1 _1491_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0709_ _0780_/A vssd1 vssd1 vccd1 vccd1 _0802_/A sky130_fd_sc_hd__inv_2
XFILLER_0_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0991_ hold147/X _1069_/S _1103_/B _0990_/X vssd1 vssd1 vccd1 vccd1 _0991_/X sky130_fd_sc_hd__a22o_1
XANTENNA__0980__A1_N _0971_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1474_ _1580_/CLK _1474_/D _1256_/Y vssd1 vssd1 vccd1 vccd1 _1474_/Q sky130_fd_sc_hd__dfrtp_1
X_1543_ _1544_/CLK _1543_/D _1325_/Y vssd1 vssd1 vccd1 vccd1 _1543_/Q sky130_fd_sc_hd__dfrtp_1
X_1612_ _1612_/CLK _1612_/D _1394_/Y vssd1 vssd1 vccd1 vccd1 _1612_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold241 _1460_/Q vssd1 vssd1 vccd1 vccd1 hold241/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 hold385/X vssd1 vssd1 vccd1 vccd1 hold263/X sky130_fd_sc_hd__buf_1
Xhold285 _0842_/X vssd1 vssd1 vccd1 vccd1 _1610_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 _1620_/Q vssd1 vssd1 vccd1 vccd1 _0813_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold274 _1618_/Q vssd1 vssd1 vccd1 vccd1 _0817_/A sky130_fd_sc_hd__buf_1
Xhold230 _1540_/Q vssd1 vssd1 vccd1 vccd1 hold230/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 _1503_/Q vssd1 vssd1 vccd1 vccd1 _1136_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput9 wb_dat_i[13] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1190_ _1192_/D _1192_/B _1192_/C _1590_/Q vssd1 vssd1 vccd1 vccd1 _1191_/C sky130_fd_sc_hd__or4b_1
XFILLER_0_54_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0974_ _0971_/Y _1015_/A hold44/X _1059_/A2 vssd1 vssd1 vccd1 vccd1 _1559_/D sky130_fd_sc_hd__a2bb2o_1
X_1457_ _1583_/CLK _1457_/D _1239_/Y vssd1 vssd1 vccd1 vccd1 _1457_/Q sky130_fd_sc_hd__dfrtp_1
X_1526_ _1547_/CLK hold87/X _1308_/Y vssd1 vssd1 vccd1 vccd1 hold42/A sky130_fd_sc_hd__dfrtp_1
X_1388_ _1409_/A vssd1 vssd1 vccd1 vccd1 _1388_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_37_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_13_clk_A clkbuf_1_1__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1068__A0 hold84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1311_ _1404_/A vssd1 vssd1 vccd1 vccd1 _1311_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_11_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1242_ _1397_/A vssd1 vssd1 vccd1 vccd1 _1242_/Y sky130_fd_sc_hd__inv_2
X_1173_ hold74/X hold102/X _1173_/S vssd1 vssd1 vccd1 vccd1 _1173_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_27_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1031__C _1031_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0888_ _0918_/C vssd1 vssd1 vccd1 vccd1 _0917_/B sky130_fd_sc_hd__inv_2
XFILLER_0_42_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout117_A _1007_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0957_ _1100_/A hold86/X _1100_/B _1100_/C vssd1 vssd1 vccd1 vccd1 _1178_/S sky130_fd_sc_hd__and4bb_2
X_1509_ _1612_/CLK _1509_/D _1291_/Y vssd1 vssd1 vccd1 vccd1 _1509_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_26_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _1558_/CLK sky130_fd_sc_hd__clkbuf_16
Xinput23 wb_dat_i[26] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__buf_1
Xinput12 wb_dat_i[16] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__clkbuf_1
X_0742_ hold54/X _0726_/A _0753_/D hold139/X vssd1 vssd1 vccd1 vccd1 _0742_/X sky130_fd_sc_hd__o31a_1
X_0811_ _0806_/A _0836_/A _0805_/Y _0776_/A vssd1 vssd1 vccd1 vccd1 _0812_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_24_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput34 wb_dat_i[7] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__buf_1
X_1225_ _1417_/A vssd1 vssd1 vccd1 vccd1 _1225_/Y sky130_fd_sc_hd__inv_2
X_1156_ hold18/X _1441_/Q _1173_/S vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_17_clk clkbuf_1_1__f_clk/X vssd1 vssd1 vccd1 vccd1 _1627_/CLK sky130_fd_sc_hd__clkbuf_16
X_1087_ _1086_/X hold141/X _1099_/S vssd1 vssd1 vccd1 vccd1 _1087_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1010_ _1100_/A hold94/X _1192_/C vssd1 vssd1 vccd1 vccd1 _1011_/B sky130_fd_sc_hd__and3b_1
XFILLER_0_56_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_6_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _1583_/CLK sky130_fd_sc_hd__clkbuf_16
X_0725_ _0882_/A hold54/X vssd1 vssd1 vccd1 vccd1 _0764_/C sky130_fd_sc_hd__or2_1
XFILLER_0_12_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1208_ _1397_/A vssd1 vssd1 vccd1 vccd1 _1208_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_18_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1139_ _1138_/A _1138_/B _1184_/A vssd1 vssd1 vccd1 vccd1 _1141_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1490_ _1602_/CLK hold61/X _1272_/Y vssd1 vssd1 vccd1 vccd1 hold60/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__0977__A _1100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1611_ _1615_/CLK _1611_/D _1393_/Y vssd1 vssd1 vccd1 vccd1 _1611_/Q sky130_fd_sc_hd__dfrtp_1
X_0990_ hold81/X _0990_/B vssd1 vssd1 vccd1 vccd1 _0990_/X sky130_fd_sc_hd__and2_1
X_1473_ _1582_/CLK _1473_/D _1255_/Y vssd1 vssd1 vccd1 vccd1 _1473_/Q sky130_fd_sc_hd__dfrtp_1
X_1542_ _1612_/CLK _1542_/D _1324_/Y vssd1 vssd1 vccd1 vccd1 _1542_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold231 _1541_/Q vssd1 vssd1 vccd1 vccd1 hold231/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 hold383/X vssd1 vssd1 vccd1 vccd1 hold253/X sky130_fd_sc_hd__buf_1
Xhold242 _1499_/Q vssd1 vssd1 vccd1 vccd1 _1137_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold220 _1549_/Q vssd1 vssd1 vccd1 vccd1 hold220/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold264 _1149_/X vssd1 vssd1 vccd1 vccd1 _1448_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold297 _0814_/X vssd1 vssd1 vccd1 vccd1 _1620_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 _0821_/X vssd1 vssd1 vccd1 vccd1 _1618_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold286 _1514_/Q vssd1 vssd1 vccd1 vccd1 hold286/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_55_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1416__A _1416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0990__A hold81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0973_ _1100_/A _1100_/C _1191_/B vssd1 vssd1 vccd1 vccd1 _1015_/A sky130_fd_sc_hd__or3b_2
XFILLER_0_10_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1525_ _1612_/CLK _1525_/D _1307_/Y vssd1 vssd1 vccd1 vccd1 hold50/A sky130_fd_sc_hd__dfrtp_1
X_1456_ _1548_/CLK _1456_/D _1238_/Y vssd1 vssd1 vccd1 vccd1 _1456_/Q sky130_fd_sc_hd__dfrtp_1
X_1387_ _1387_/A vssd1 vssd1 vccd1 vccd1 _1387_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_26_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1310_ _1404_/A vssd1 vssd1 vccd1 vccd1 _1310_/Y sky130_fd_sc_hd__inv_2
X_1241_ _1387_/A vssd1 vssd1 vccd1 vccd1 _1241_/Y sky130_fd_sc_hd__inv_2
XANTENNA__0985__A _1100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1059__B2 hold165/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1172_ hold92/X hold151/X _1173_/S vssd1 vssd1 vccd1 vccd1 _1172_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_42_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0956_ _1100_/A _0954_/Y _0955_/X vssd1 vssd1 vccd1 vccd1 _1564_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_12_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput100 _1463_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[7] sky130_fd_sc_hd__buf_12
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0887_ _0889_/C _0887_/B _0915_/C vssd1 vssd1 vccd1 vccd1 _0918_/C sky130_fd_sc_hd__and3_1
XFILLER_0_2_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1439_ _1634_/CLK _1439_/D _1221_/Y vssd1 vssd1 vccd1 vccd1 _1439_/Q sky130_fd_sc_hd__dfrtp_1
X_1508_ _1558_/CLK _1508_/D _1290_/Y vssd1 vssd1 vccd1 vccd1 hold88/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput13 wb_dat_i[17] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_56_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0810_ _0810_/A _0810_/B vssd1 vssd1 vccd1 vccd1 _0810_/X sky130_fd_sc_hd__and2_1
XANTENNA__0971__C _1103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0741_ _0917_/A _0741_/B _0741_/C _0906_/B vssd1 vssd1 vccd1 vccd1 _0764_/D sky130_fd_sc_hd__or4_1
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput24 wb_dat_i[27] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__clkbuf_1
Xinput35 wb_dat_i[8] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__buf_1
XFILLER_0_42_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1224_ _1409_/A vssd1 vssd1 vccd1 vccd1 _1224_/Y sky130_fd_sc_hd__inv_2
X_1155_ hold232/X _1442_/Q _1168_/S vssd1 vssd1 vccd1 vccd1 _1155_/X sky130_fd_sc_hd__mux2_1
X_1086_ _1098_/A _1086_/B vssd1 vssd1 vccd1 vccd1 _1086_/X sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_12_clk_A clkbuf_1_1__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0939_ _0967_/B _1141_/A vssd1 vssd1 vccd1 vccd1 _0939_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_2_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_27_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0724_ _0764_/A _0884_/S vssd1 vssd1 vccd1 vccd1 _0726_/A sky130_fd_sc_hd__or2_2
XFILLER_0_8_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1207_ _1417_/A vssd1 vssd1 vccd1 vccd1 _1207_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_18_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1069_ hold371/X _1137_/B _1069_/S vssd1 vssd1 vccd1 vccd1 _1069_/X sky130_fd_sc_hd__mux2_1
X_1138_ _1138_/A _1138_/B vssd1 vssd1 vccd1 vccd1 _1184_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_47_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0977__B _1007_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1181__B1_N _1173_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0993__A hold81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1610_ _1623_/CLK _1610_/D _1392_/Y vssd1 vssd1 vccd1 vccd1 _1610_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1541_ _1612_/CLK _1541_/D _1323_/Y vssd1 vssd1 vccd1 vccd1 _1541_/Q sky130_fd_sc_hd__dfrtp_1
X_1472_ _1601_/CLK hold11/X _1254_/Y vssd1 vssd1 vccd1 vccd1 _1472_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0992__A_N _1100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold254 _1144_/X vssd1 vssd1 vccd1 vccd1 _1453_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 hold376/X vssd1 vssd1 vccd1 vccd1 hold265/X sky130_fd_sc_hd__buf_1
XFILLER_0_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold210 _1629_/Q vssd1 vssd1 vccd1 vccd1 hold210/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 _1523_/Q vssd1 vssd1 vccd1 vccd1 hold232/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold243 _1069_/X vssd1 vssd1 vccd1 vccd1 _1499_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 _1627_/Q vssd1 vssd1 vccd1 vccd1 _0847_/A sky130_fd_sc_hd__clkbuf_2
Xhold287 _1164_/X vssd1 vssd1 vccd1 vccd1 _1433_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 _1420_/Q vssd1 vssd1 vccd1 vccd1 _1141_/A sky130_fd_sc_hd__clkbuf_2
Xhold298 _1582_/Q vssd1 vssd1 vccd1 vccd1 _0739_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0972_ _1013_/A _0971_/Y hold175/X _1061_/A2 vssd1 vssd1 vccd1 vccd1 _1560_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_6_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1524_ _1586_/CLK _1524_/D _1306_/Y vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1455_ _1558_/CLK _1455_/D _1237_/Y vssd1 vssd1 vccd1 vccd1 _1455_/Q sky130_fd_sc_hd__dfrtp_1
X_1386_ _1409_/A vssd1 vssd1 vccd1 vccd1 _1386_/Y sky130_fd_sc_hd__inv_2
XANTENNA__0976__A2_N _0975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0969__C _1007_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1171_ hold68/X _1426_/Q _1171_/S vssd1 vssd1 vccd1 vccd1 hold69/A sky130_fd_sc_hd__mux2_1
X_1240_ _1387_/A vssd1 vssd1 vccd1 vccd1 _1240_/Y sky130_fd_sc_hd__inv_2
XANTENNA__0985__B _1100_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1059__A2 _1059_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0886_ _0886_/A _0886_/B _0886_/C _0935_/S vssd1 vssd1 vccd1 vccd1 _0915_/C sky130_fd_sc_hd__and4_2
XFILLER_0_6_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0955_ _1100_/A _0966_/S _0955_/C _0963_/B vssd1 vssd1 vccd1 vccd1 _0955_/X sky130_fd_sc_hd__and4b_1
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1507_ _1544_/CLK _1507_/D _1289_/Y vssd1 vssd1 vccd1 vccd1 hold68/A sky130_fd_sc_hd__dfrtp_1
Xoutput101 _1464_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[8] sky130_fd_sc_hd__buf_12
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1438_ _1583_/CLK _1438_/D _1220_/Y vssd1 vssd1 vccd1 vccd1 _1438_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1369_ _1413_/A vssd1 vssd1 vccd1 vccd1 _1369_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput14 wb_dat_i[18] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0740_ _0740_/A _0740_/B _0740_/C _0740_/D vssd1 vssd1 vccd1 vccd1 _0906_/B sky130_fd_sc_hd__or4_1
XFILLER_0_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput36 wb_dat_i[9] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__clkbuf_1
Xinput25 wb_dat_i[28] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__buf_1
XANTENNA__0996__A hold81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1154_ hold28/X _1443_/Q _1173_/S vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__mux2_1
X_1223_ _1415_/A vssd1 vssd1 vccd1 vccd1 _1223_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_23_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1085_ input31/X input8/X input17/X input25/X _1100_/C _1100_/B vssd1 vssd1 vccd1
+ vccd1 _1086_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_30_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout122_A _1416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0869_ _1592_/Q hold2/X _0874_/S vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__mux2_1
XFILLER_0_23_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0938_ _1488_/Q _1101_/B vssd1 vssd1 vccd1 vccd1 _0938_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_38_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0723_ _0764_/A _0884_/S vssd1 vssd1 vccd1 vccd1 _0882_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_8_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1137_ _1187_/D _1137_/B _1187_/C _1137_/D vssd1 vssd1 vccd1 vccd1 _1138_/B sky130_fd_sc_hd__and4b_1
X_1206_ _1339_/A vssd1 vssd1 vccd1 vccd1 _1206_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_34_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1068_ hold84/X _1187_/D _1068_/S vssd1 vssd1 vccd1 vccd1 _1500_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_11_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_11_clk_A clkbuf_1_1__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_26_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1022__B1 _1103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1540_ _1605_/CLK _1540_/D _1322_/Y vssd1 vssd1 vccd1 vccd1 _1540_/Q sky130_fd_sc_hd__dfrtp_1
X_1471_ _1505_/CLK _1471_/D _1253_/Y vssd1 vssd1 vccd1 vccd1 _1471_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1104__S _1135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold299 _0730_/X vssd1 vssd1 vccd1 vccd1 _0733_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 _1481_/Q vssd1 vssd1 vccd1 vccd1 hold288/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 _1162_/X vssd1 vssd1 vccd1 vccd1 _1435_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold255 hold378/X vssd1 vssd1 vccd1 vccd1 _1192_/B sky130_fd_sc_hd__clkbuf_2
Xhold211 _0873_/X vssd1 vssd1 vccd1 vccd1 _1588_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 _1155_/X vssd1 vssd1 vccd1 vccd1 _1442_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold222 _1200_/Y vssd1 vssd1 vccd1 vccd1 _1606_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold200 _1512_/Q vssd1 vssd1 vccd1 vccd1 hold200/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold244 _1502_/Q vssd1 vssd1 vccd1 vccd1 _1188_/C sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1075__A _1100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold277 _1029_/B vssd1 vssd1 vccd1 vccd1 hold277/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0971_ hold86/X hold80/X _1103_/B vssd1 vssd1 vccd1 vccd1 _0971_/Y sky130_fd_sc_hd__nand3b_4
X_1523_ _1598_/CLK _1523_/D _1305_/Y vssd1 vssd1 vccd1 vccd1 _1523_/Q sky130_fd_sc_hd__dfrtp_1
X_1454_ _1556_/CLK _1454_/D _1236_/Y vssd1 vssd1 vccd1 vccd1 _1454_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__0999__A hold81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1385_ _1385_/A vssd1 vssd1 vccd1 vccd1 _1385_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_45_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1170_ hold88/X _1427_/Q _1173_/S vssd1 vssd1 vccd1 vccd1 hold89/A sky130_fd_sc_hd__mux2_1
X_0885_ _0886_/B _1568_/Q _1567_/Q vssd1 vssd1 vccd1 vccd1 _0885_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_2_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0954_ _0955_/C _0953_/Y _0966_/S vssd1 vssd1 vccd1 vccd1 _0954_/Y sky130_fd_sc_hd__o21ai_1
X_1437_ _1612_/CLK hold47/X _1219_/Y vssd1 vssd1 vccd1 vccd1 _1437_/Q sky130_fd_sc_hd__dfrtp_1
X_1506_ _1586_/CLK hold93/X _1288_/Y vssd1 vssd1 vccd1 vccd1 hold92/A sky130_fd_sc_hd__dfrtp_1
Xoutput102 hold96/A vssd1 vssd1 vccd1 vccd1 wb_dat_o[9] sky130_fd_sc_hd__buf_12
X_1368_ _1417_/A vssd1 vssd1 vccd1 vccd1 _1368_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_37_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1299_ _1339_/A vssd1 vssd1 vccd1 vccd1 _1299_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_18_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput15 wb_dat_i[19] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput26 wb_dat_i[29] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1010__A_N _1100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1153_ hold50/X _1444_/Q _1168_/S vssd1 vssd1 vccd1 vccd1 hold51/A sky130_fd_sc_hd__mux2_1
X_1222_ _1385_/A vssd1 vssd1 vccd1 vccd1 _1222_/Y sky130_fd_sc_hd__inv_2
X_1084_ _1083_/X hold104/X _1096_/S vssd1 vssd1 vccd1 vccd1 _1084_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1112__S _1135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_9_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _1589_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_30_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0799_ _0803_/D _0837_/A _0837_/B _0804_/C vssd1 vssd1 vccd1 vccd1 _0817_/D sky130_fd_sc_hd__and4_1
X_0868_ _1593_/Q hold4/X _0874_/S vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__mux2_1
XFILLER_0_2_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0937_ hold346/X _0967_/B _1141_/A vssd1 vssd1 vccd1 vccd1 _1101_/C sky130_fd_sc_hd__and3b_2
XFILLER_0_38_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0722_ _1387_/A vssd1 vssd1 vccd1 vccd1 _0722_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_12_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1107__S _1133_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1205_ _1402_/A vssd1 vssd1 vccd1 vccd1 _1205_/Y sky130_fd_sc_hd__inv_2
X_1067_ _1192_/D _1136_/D _1071_/S vssd1 vssd1 vccd1 vccd1 _1501_/D sky130_fd_sc_hd__mux2_1
X_1136_ _1188_/D _1136_/B _1188_/C _1136_/D vssd1 vssd1 vccd1 vccd1 _1138_/A sky130_fd_sc_hd__and4b_1
XFILLER_0_50_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1119_ hold10/X _1472_/Q _1133_/S vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__mux2_1
XFILLER_0_41_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1470_ _1634_/CLK hold77/X _1252_/Y vssd1 vssd1 vccd1 vccd1 _1470_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold201 _1056_/X vssd1 vssd1 vccd1 vccd1 _1512_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1120__S _1133_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold245 _1578_/Q vssd1 vssd1 vccd1 vccd1 _0892_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold289 _1576_/Q vssd1 vssd1 vccd1 vccd1 _0914_/S sky130_fd_sc_hd__buf_1
Xhold212 _1555_/Q vssd1 vssd1 vccd1 vccd1 hold212/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 _1572_/Q vssd1 vssd1 vccd1 vccd1 _0889_/C sky130_fd_sc_hd__buf_1
Xhold256 _1488_/Q vssd1 vssd1 vccd1 vccd1 _0775_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 _1626_/Q vssd1 vssd1 vccd1 vccd1 _0850_/A sky130_fd_sc_hd__clkbuf_2
Xhold234 _1536_/Q vssd1 vssd1 vccd1 vccd1 hold234/X sky130_fd_sc_hd__dlygate4sd3_1
X_1599_ _1624_/CLK hold33/X _1381_/Y vssd1 vssd1 vccd1 vccd1 hold32/A sky130_fd_sc_hd__dfrtp_1
Xhold223 _1501_/Q vssd1 vssd1 vccd1 vccd1 _1136_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_56_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0975__C_N _0995_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_10_clk_A clkbuf_1_1__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_25_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0970_ _1140_/A _1185_/B vssd1 vssd1 vccd1 vccd1 _0970_/X sky130_fd_sc_hd__and2_2
X_1453_ _1612_/CLK _1453_/D _1235_/Y vssd1 vssd1 vccd1 vccd1 _1453_/Q sky130_fd_sc_hd__dfrtp_1
X_1522_ _1586_/CLK _1522_/D _1304_/Y vssd1 vssd1 vccd1 vccd1 _1522_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1115__S _1133_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1384_ _1384_/A vssd1 vssd1 vccd1 vccd1 _1384_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_42_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput103 _1636_/X vssd1 vssd1 vccd1 vccd1 wb_stb_o sky130_fd_sc_hd__buf_12
XFILLER_0_42_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0884_ _0735_/Y _0880_/B _0884_/S vssd1 vssd1 vccd1 vccd1 _1583_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_2_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0953_ _0963_/B vssd1 vssd1 vccd1 vccd1 _0953_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_10_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1367_ _1417_/A vssd1 vssd1 vccd1 vccd1 _1367_/Y sky130_fd_sc_hd__inv_2
X_1505_ _1505_/CLK hold75/X _1287_/Y vssd1 vssd1 vccd1 vccd1 hold74/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1436_ _1556_/CLK hold35/X _1218_/Y vssd1 vssd1 vccd1 vccd1 _1436_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1298_ _1413_/A vssd1 vssd1 vccd1 vccd1 _1298_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_33_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0966__A0 _1007_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput16 wb_dat_i[1] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__buf_1
Xinput27 wb_dat_i[2] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1221_ _1415_/A vssd1 vssd1 vccd1 vccd1 _1221_/Y sky130_fd_sc_hd__inv_2
X_1152_ hold42/X _1445_/Q _1168_/S vssd1 vssd1 vccd1 vccd1 hold43/A sky130_fd_sc_hd__mux2_1
X_1083_ _1098_/A _1083_/B vssd1 vssd1 vccd1 vccd1 _1083_/X sky130_fd_sc_hd__and2_1
X_0936_ _0936_/A vssd1 vssd1 vccd1 vccd1 _1567_/D sky130_fd_sc_hd__inv_2
XFILLER_0_23_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0798_ _0828_/A _0833_/A _0798_/C vssd1 vssd1 vccd1 vccd1 _0804_/C sky130_fd_sc_hd__and3_1
X_0867_ hold367/X hold139/X _0874_/S vssd1 vssd1 vccd1 vccd1 _0867_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_30_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout108_A _1129_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1419_ _1489_/CLK _1419_/D _1201_/Y vssd1 vssd1 vccd1 vccd1 _1419_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0721_ _0933_/B vssd1 vssd1 vccd1 vccd1 _0917_/A sky130_fd_sc_hd__inv_2
XFILLER_0_12_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1204_ _1410_/A vssd1 vssd1 vccd1 vccd1 _1204_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_18_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1135_ hold112/X hold133/X _1135_/S vssd1 vssd1 vccd1 vccd1 _1135_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1123__S _1133_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1066_ _0995_/C _1188_/C _1071_/S vssd1 vssd1 vccd1 vccd1 _1502_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_50_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0919_ _0919_/A _0919_/B vssd1 vssd1 vccd1 vccd1 _0919_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_7_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0974__A2_N _1015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1118__S _1135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1118_ hold225/X _1473_/Q _1135_/S vssd1 vssd1 vccd1 vccd1 _1118_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_35_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1049_ hold202/X _1069_/S hold82/X _1031_/C vssd1 vssd1 vccd1 vccd1 _1519_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_43_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1022__A2 _1069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold213 _1117_/X vssd1 vssd1 vccd1 vccd1 _1474_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold202 _1519_/Q vssd1 vssd1 vccd1 vccd1 hold202/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold224 _1468_/Q vssd1 vssd1 vccd1 vccd1 hold224/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 _1142_/X vssd1 vssd1 vccd1 vccd1 _1455_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 _0909_/X vssd1 vssd1 vccd1 vccd1 _1578_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 _0926_/X vssd1 vssd1 vccd1 vccd1 _1572_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1598_ _1598_/CLK _1598_/D _1380_/Y vssd1 vssd1 vccd1 vccd1 _1598_/Q sky130_fd_sc_hd__dfrtp_1
Xhold279 _0850_/X vssd1 vssd1 vccd1 vccd1 _0852_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 _1102_/X vssd1 vssd1 vccd1 vccd1 _1488_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1521_ _1600_/CLK _1521_/D _1303_/Y vssd1 vssd1 vccd1 vccd1 _1521_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1452_ _1562_/CLK hold99/X _1234_/Y vssd1 vssd1 vccd1 vccd1 _1452_/Q sky130_fd_sc_hd__dfrtp_1
X_1383_ _1384_/A vssd1 vssd1 vccd1 vccd1 _1383_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1131__S _1135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0984__B2 _1071_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0952_ _1101_/C _1185_/B _1029_/B vssd1 vssd1 vccd1 vccd1 _0963_/B sky130_fd_sc_hd__or3_2
XFILLER_0_50_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0883_ _0764_/A _0880_/B _0882_/X vssd1 vssd1 vccd1 vccd1 _1584_/D sky130_fd_sc_hd__a21bo_1
Xoutput104 _1423_/Q vssd1 vssd1 vccd1 vccd1 wb_we_o sky130_fd_sc_hd__buf_12
X_1504_ _1632_/CLK _1504_/D _1286_/Y vssd1 vssd1 vccd1 vccd1 _1504_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1435_ _1586_/CLK _1435_/D _1217_/Y vssd1 vssd1 vccd1 vccd1 _1435_/Q sky130_fd_sc_hd__dfrtp_1
X_1366_ _1417_/A vssd1 vssd1 vccd1 vccd1 _1366_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_37_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1126__S _1133_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1297_ _1405_/A vssd1 vssd1 vccd1 vccd1 _1297_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_33_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_24_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput17 wb_dat_i[20] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__buf_1
XFILLER_0_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput28 wb_dat_i[30] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__buf_1
X_1220_ _1417_/A vssd1 vssd1 vccd1 vccd1 _1220_/Y sky130_fd_sc_hd__inv_2
X_1151_ hold70/X _1446_/Q _1168_/S vssd1 vssd1 vccd1 vccd1 hold71/A sky130_fd_sc_hd__mux2_1
X_1082_ input32/X input9/X input18/X input26/X _1100_/C _1100_/B vssd1 vssd1 vccd1
+ vccd1 _1083_/B sky130_fd_sc_hd__mux4_1
X_0935_ _0925_/A _0933_/B _0935_/S vssd1 vssd1 vccd1 vccd1 _0936_/A sky130_fd_sc_hd__mux2_1
X_0866_ _0866_/A _0882_/C vssd1 vssd1 vccd1 vccd1 _0874_/S sky130_fd_sc_hd__nor2_4
XANTENNA__1070__A0 _1007_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0797_ _0837_/A _0837_/B vssd1 vssd1 vccd1 vccd1 _0831_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_30_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1349_ _1363_/A vssd1 vssd1 vccd1 vccd1 _1349_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_48_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1418_ _1632_/CLK _1418_/D _0722_/Y vssd1 vssd1 vccd1 vccd1 _1418_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1061__B1 _1023_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0720_ input4/X vssd1 vssd1 vccd1 vccd1 _0720_/Y sky130_fd_sc_hd__inv_2
XANTENNA_output99_A _1462_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1134_ hold149/X hold181/X _1135_/S vssd1 vssd1 vccd1 vccd1 _1134_/X sky130_fd_sc_hd__mux2_1
X_1203_ _1402_/A vssd1 vssd1 vccd1 vccd1 _1203_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1065_ _1191_/B _1136_/B _1071_/S vssd1 vssd1 vccd1 vccd1 _1503_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_55_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0918_ _0923_/S _0933_/B _0918_/C vssd1 vssd1 vccd1 vccd1 _0920_/S sky130_fd_sc_hd__and3_1
XANTENNA_fanout120_A _1416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0849_ _0789_/A _0849_/B vssd1 vssd1 vccd1 vccd1 _0855_/A sky130_fd_sc_hd__and2b_1
XANTENNA_hold165_A _1029_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_10_clk clkbuf_1_1__f_clk/X vssd1 vssd1 vccd1 vccd1 _1548_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1117_ hold212/X _1474_/Q _1135_/S vssd1 vssd1 vccd1 vccd1 _1117_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1134__S _1135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1016__B1 _0970_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1048_ hold100/X _1069_/S _0990_/X _1031_/C vssd1 vssd1 vccd1 vccd1 _1048_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_1__f_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_26_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold247 _1580_/Q vssd1 vssd1 vccd1 vccd1 _0893_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold203 _1159_/X vssd1 vssd1 vccd1 vccd1 _1438_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1129__S _1129_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold225 _1554_/Q vssd1 vssd1 vccd1 vccd1 hold225/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold269 _1487_/Q vssd1 vssd1 vccd1 vccd1 hold269/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 _1500_/Q vssd1 vssd1 vccd1 vccd1 _1187_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold236 _1535_/Q vssd1 vssd1 vccd1 vccd1 hold236/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 _1492_/Q vssd1 vssd1 vccd1 vccd1 hold214/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1597_ _1602_/CLK hold49/X _1379_/Y vssd1 vssd1 vccd1 vccd1 hold48/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1520_ _1556_/CLK _1520_/D _1302_/Y vssd1 vssd1 vccd1 vccd1 _1520_/Q sky130_fd_sc_hd__dfrtp_1
X_1451_ _1548_/CLK hold79/X _1233_/Y vssd1 vssd1 vccd1 vccd1 hold78/A sky130_fd_sc_hd__dfrtp_2
X_1382_ _1384_/A vssd1 vssd1 vccd1 vccd1 _1382_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_45_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0882_ _0882_/A _0882_/B _0882_/C _0880_/A vssd1 vssd1 vccd1 vccd1 _0882_/X sky130_fd_sc_hd__or4b_1
X_0951_ _1420_/Q _1418_/Q hold363/X vssd1 vssd1 vccd1 vccd1 _1184_/A sky130_fd_sc_hd__or3b_1
XFILLER_0_2_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1503_ _1632_/CLK _1503_/D _1285_/Y vssd1 vssd1 vccd1 vccd1 _1503_/Q sky130_fd_sc_hd__dfrtp_1
X_1434_ _1544_/CLK _1434_/D _1216_/Y vssd1 vssd1 vccd1 vccd1 _1434_/Q sky130_fd_sc_hd__dfrtp_1
X_1365_ _1417_/A vssd1 vssd1 vccd1 vccd1 _1365_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_37_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1296_ _1415_/A vssd1 vssd1 vccd1 vccd1 _1296_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1142__S _1173_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 wb_dat_i[21] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__buf_1
XFILLER_0_32_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput29 wb_dat_i[31] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__buf_1
X_1150_ hold239/X _1447_/Q _1168_/S vssd1 vssd1 vccd1 vccd1 _1150_/X sky130_fd_sc_hd__mux2_1
X_1081_ _1080_/X hold20/X _1099_/S vssd1 vssd1 vccd1 vccd1 _1081_/X sky130_fd_sc_hd__mux2_1
X_0934_ _0886_/C _0913_/A _0933_/X _0932_/Y _0917_/A vssd1 vssd1 vccd1 vccd1 _0934_/X
+ sky130_fd_sc_hd__o32a_1
X_0865_ hold369/X hold8/X _0865_/S vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__mux2_1
XFILLER_0_23_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0796_ _0837_/B vssd1 vssd1 vccd1 vccd1 _0796_/Y sky130_fd_sc_hd__inv_2
X_1417_ _1417_/A vssd1 vssd1 vccd1 vccd1 _1417_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_2_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1348_ _1413_/A vssd1 vssd1 vccd1 vccd1 _1348_/Y sky130_fd_sc_hd__inv_2
X_1279_ _1413_/A vssd1 vssd1 vccd1 vccd1 _1279_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1061__B2 hold165/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1052__B2 _1031_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_23_clk_A clkbuf_1_1__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1133_ hold64/X hold169/X _1133_/S vssd1 vssd1 vccd1 vccd1 _1133_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_18_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1064_ _0989_/C _1188_/D _1071_/S vssd1 vssd1 vccd1 vccd1 _1504_/D sky130_fd_sc_hd__mux2_1
X_1202_ _1384_/A vssd1 vssd1 vccd1 vccd1 _1202_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1043__B2 _1059_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0917_ _0917_/A _0917_/B vssd1 vssd1 vccd1 vccd1 _0917_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_fanout113_A _1059_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0779_ _0803_/A _0817_/A _0822_/A _0803_/D vssd1 vssd1 vccd1 vccd1 _0781_/C sky130_fd_sc_hd__or4_1
X_0848_ _0851_/S _1596_/Q _0847_/Y _0846_/X _0850_/A vssd1 vssd1 vccd1 vccd1 _0849_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_38_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1034__B2 _1030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1150__S _1168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1047_ hold118/X _1031_/Y hold216/X _1059_/A2 vssd1 vssd1 vccd1 vccd1 _1521_/D sky130_fd_sc_hd__a2bb2o_1
X_1116_ hold22/X _1475_/Q _1133_/S vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__mux2_1
XANTENNA__1016__B2 _1015_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold248 _0904_/X vssd1 vssd1 vccd1 vccd1 _1580_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 _1118_/X vssd1 vssd1 vccd1 vccd1 _1473_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold259 hold381/X vssd1 vssd1 vccd1 vccd1 hold259/X sky130_fd_sc_hd__buf_1
Xhold204 _1462_/Q vssd1 vssd1 vccd1 vccd1 hold204/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1596_ _1598_/CLK hold9/X _1378_/Y vssd1 vssd1 vccd1 vccd1 _1596_/Q sky130_fd_sc_hd__dfrtp_1
Xhold237 _1459_/Q vssd1 vssd1 vccd1 vccd1 hold237/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 _1090_/X vssd1 vssd1 vccd1 vccd1 _1492_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1145__S _1173_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1450_ _1586_/CLK hold73/X _1232_/Y vssd1 vssd1 vccd1 vccd1 _1450_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1381_ _1385_/A vssd1 vssd1 vccd1 vccd1 _1381_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1164__A0 hold286/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1579_ _1582_/CLK _1579_/D _1361_/Y vssd1 vssd1 vccd1 vccd1 _1579_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0881_ hold54/X _0880_/Y hold262/X vssd1 vssd1 vccd1 vccd1 _1585_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_2_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0950_ _1141_/A _0950_/B _0967_/B vssd1 vssd1 vccd1 vccd1 _1029_/B sky130_fd_sc_hd__nor3b_1
XFILLER_0_10_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1502_ _1562_/CLK _1502_/D _1284_/Y vssd1 vssd1 vccd1 vccd1 _1502_/Q sky130_fd_sc_hd__dfrtp_1
X_1433_ _1624_/CLK _1433_/D _1215_/Y vssd1 vssd1 vccd1 vccd1 _1433_/Q sky130_fd_sc_hd__dfrtp_1
X_1364_ _1364_/A vssd1 vssd1 vccd1 vccd1 _1364_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_37_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1295_ _1409_/A vssd1 vssd1 vccd1 vccd1 _1295_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_53_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0972__A2_N _0971_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0998__A_N _1100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput19 wb_dat_i[22] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__buf_1
X_1080_ _1098_/A _1080_/B vssd1 vssd1 vccd1 vccd1 _1080_/X sky130_fd_sc_hd__and2_1
XFILLER_0_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0933_ _1567_/Q _0933_/B vssd1 vssd1 vccd1 vccd1 _0933_/X sky130_fd_sc_hd__and2_1
X_0795_ _0795_/A _0795_/B _0843_/A _0845_/S vssd1 vssd1 vccd1 vccd1 _0837_/B sky130_fd_sc_hd__and4_2
XFILLER_0_23_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0864_ hold48/X hold60/X _0865_/S vssd1 vssd1 vccd1 vccd1 hold49/A sky130_fd_sc_hd__mux2_1
X_1416_ _1416_/A vssd1 vssd1 vccd1 vccd1 _1416_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_23_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1347_ _1385_/A vssd1 vssd1 vccd1 vccd1 _1347_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1153__S _1168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1278_ _1385_/A vssd1 vssd1 vccd1 vccd1 _1278_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout130 _1416_/A vssd1 vssd1 vccd1 vccd1 _1409_/A sky130_fd_sc_hd__buf_6
XFILLER_0_49_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1052__A2 _1071_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1201_ _1384_/A vssd1 vssd1 vccd1 vccd1 _1201_/Y sky130_fd_sc_hd__inv_2
X_1132_ hold230/X hold237/X _1135_/S vssd1 vssd1 vccd1 vccd1 _1459_/D sky130_fd_sc_hd__mux2_1
X_1063_ hold74/X _1069_/S _1027_/Y _1031_/C vssd1 vssd1 vccd1 vccd1 hold75/A sky130_fd_sc_hd__a22o_1
XFILLER_0_18_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0916_ _0912_/A _0913_/Y _0915_/X vssd1 vssd1 vccd1 vccd1 _0916_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_50_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1002__A hold81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1148__S _1173_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0778_ _0795_/A _0843_/A _1608_/Q _0795_/B vssd1 vssd1 vccd1 vccd1 _0781_/B sky130_fd_sc_hd__or4bb_1
XANTENNA_fanout106_A _1171_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0847_ _0847_/A _0850_/A vssd1 vssd1 vccd1 vccd1 _0847_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_38_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_37_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1042__A1_N _0975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1046_ _1025_/A _1031_/Y hold18/X _1071_/S vssd1 vssd1 vccd1 vccd1 _1522_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_0_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1115_ hold38/X _1476_/Q _1133_/S vssd1 vssd1 vccd1 vccd1 hold39/A sky130_fd_sc_hd__mux2_1
XFILLER_0_43_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_22_clk_A clkbuf_1_1__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold205 _1129_/X vssd1 vssd1 vccd1 vccd1 _1462_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold249 _1498_/Q vssd1 vssd1 vccd1 vccd1 _1187_/C sky130_fd_sc_hd__dlygate4sd3_1
X_1595_ _1632_/CLK _1595_/D _1377_/Y vssd1 vssd1 vccd1 vccd1 _1595_/Q sky130_fd_sc_hd__dfrtp_1
Xhold227 _1619_/Q vssd1 vssd1 vccd1 vccd1 _0803_/A sky130_fd_sc_hd__buf_1
Xhold238 _1504_/Q vssd1 vssd1 vccd1 vccd1 _1188_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold216 _1521_/Q vssd1 vssd1 vccd1 vccd1 hold216/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_56_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1161__S _1173_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1029_ _1140_/A _1029_/B vssd1 vssd1 vccd1 vccd1 _1029_/X sky130_fd_sc_hd__and2_2
XFILLER_0_31_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1071__S _1071_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1100__A _1100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1380_ _1402_/A vssd1 vssd1 vccd1 vccd1 _1380_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0978__B2 _1069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1578_ _1580_/CLK _1578_/D _1360_/Y vssd1 vssd1 vccd1 vccd1 _1578_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1156__S _1173_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1091__A0 input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1066__S _1071_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0880_ _0880_/A _0880_/B vssd1 vssd1 vccd1 vccd1 _0880_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_27_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1363_ _1363_/A vssd1 vssd1 vccd1 vccd1 _1363_/Y sky130_fd_sc_hd__inv_2
X_1432_ _1627_/CLK _1432_/D _1214_/Y vssd1 vssd1 vccd1 vccd1 _1432_/Q sky130_fd_sc_hd__dfrtp_1
X_1501_ _1562_/CLK _1501_/D _1283_/Y vssd1 vssd1 vccd1 vccd1 _1501_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1005__A hold81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1294_ _1384_/A vssd1 vssd1 vccd1 vccd1 _1294_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_33_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0932_ _0886_/C _1567_/Q _0906_/B vssd1 vssd1 vccd1 vccd1 _0932_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_23_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0794_ _0795_/B _1609_/Q _1608_/Q vssd1 vssd1 vccd1 vccd1 _0794_/Y sky130_fd_sc_hd__nand3_1
X_0863_ hold368/X hold135/X _0865_/S vssd1 vssd1 vccd1 vccd1 _0863_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1415_ _1415_/A vssd1 vssd1 vccd1 vccd1 _1415_/Y sky130_fd_sc_hd__inv_2
X_1346_ _1387_/A vssd1 vssd1 vccd1 vccd1 _1346_/Y sky130_fd_sc_hd__inv_2
X_1277_ _1384_/A vssd1 vssd1 vccd1 vccd1 _1277_/Y sky130_fd_sc_hd__inv_2
Xfanout131 _1405_/A vssd1 vssd1 vccd1 vccd1 _1404_/A sky130_fd_sc_hd__buf_6
Xfanout120 _1416_/A vssd1 vssd1 vccd1 vccd1 _1415_/A sky130_fd_sc_hd__buf_8
XFILLER_0_14_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_22_clk clkbuf_1_1__f_clk/X vssd1 vssd1 vccd1 vccd1 _1602_/CLK sky130_fd_sc_hd__clkbuf_16
X_1200_ _0847_/A _0784_/B _0850_/X _0831_/A vssd1 vssd1 vccd1 vccd1 _1200_/Y sky130_fd_sc_hd__a31oi_1
X_1131_ hold231/X hold241/X _1135_/S vssd1 vssd1 vccd1 vccd1 _1460_/D sky130_fd_sc_hd__mux2_1
X_1062_ hold92/X _1068_/S _1025_/Y _1031_/C vssd1 vssd1 vccd1 vccd1 hold93/A sky130_fd_sc_hd__a22o_1
XFILLER_0_55_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0915_ _0912_/A _0933_/B _0915_/C _0915_/D vssd1 vssd1 vccd1 vccd1 _0915_/X sky130_fd_sc_hd__and4b_1
XANTENNA__1028__B1 _1103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_13_clk clkbuf_1_1__f_clk/X vssd1 vssd1 vccd1 vccd1 _1615_/CLK sky130_fd_sc_hd__clkbuf_16
X_0777_ _0828_/A _0835_/A _0837_/A _0833_/A vssd1 vssd1 vccd1 vccd1 _0781_/A sky130_fd_sc_hd__or4b_1
X_0846_ hold32/X hold124/X _0851_/S vssd1 vssd1 vccd1 vccd1 _0846_/X sky130_fd_sc_hd__mux2_1
X_1329_ _1385_/A vssd1 vssd1 vccd1 vccd1 _1329_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1164__S _1168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_2_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _1632_/CLK sky130_fd_sc_hd__clkbuf_16
X_1114_ hold66/X _1477_/Q _1133_/S vssd1 vssd1 vccd1 vccd1 hold67/A sky130_fd_sc_hd__mux2_1
X_1045_ _1023_/A _1031_/Y hold232/X _1061_/A2 vssd1 vssd1 vccd1 vccd1 _1523_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_0_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1159__S _1173_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0829_ _0828_/Y _0828_/A _0829_/S vssd1 vssd1 vccd1 vccd1 _0829_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_28_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1069__S _1069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold206 _1428_/Q vssd1 vssd1 vccd1 vccd1 hold206/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold217 _1157_/X vssd1 vssd1 vccd1 vccd1 _1440_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold239 _1528_/Q vssd1 vssd1 vccd1 vccd1 hold239/X sky130_fd_sc_hd__dlygate4sd3_1
X_1594_ _1635_/CLK _1594_/D _1376_/Y vssd1 vssd1 vccd1 vccd1 _1594_/Q sky130_fd_sc_hd__dfrtp_1
Xhold228 _0819_/Y vssd1 vssd1 vccd1 vccd1 _1619_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1008__A hold81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1028_ hold112/X _1061_/A2 _1103_/B _1027_/Y vssd1 vssd1 vccd1 vccd1 _1028_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1041__A1_N _1015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1100__B _1100_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1577_ _1580_/CLK _1577_/D _1359_/Y vssd1 vssd1 vccd1 vccd1 _1577_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1172__S _1173_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_21_clk_A clkbuf_1_1__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1082__A1 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1500_ _1632_/CLK _1500_/D _1282_/Y vssd1 vssd1 vccd1 vccd1 _1500_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1362_ _1364_/A vssd1 vssd1 vccd1 vccd1 _1362_/Y sky130_fd_sc_hd__inv_2
Xoutput90 _1483_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[27] sky130_fd_sc_hd__buf_12
X_1431_ _1601_/CLK _1431_/D _1213_/Y vssd1 vssd1 vccd1 vccd1 _1431_/Q sky130_fd_sc_hd__dfrtp_1
X_1293_ _1385_/A vssd1 vssd1 vccd1 vccd1 _1293_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_53_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1629_ _1631_/CLK _1629_/D _1411_/Y vssd1 vssd1 vccd1 vccd1 _1629_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1167__S _1168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0931_ _0885_/Y _0906_/X _0930_/X _0925_/A _0886_/B vssd1 vssd1 vccd1 vccd1 _0931_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__1055__B2 _1031_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0862_ hold32/X hold214/X _0865_/S vssd1 vssd1 vccd1 vccd1 hold33/A sky130_fd_sc_hd__mux2_1
XFILLER_0_48_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0793_ _0843_/A _1608_/Q vssd1 vssd1 vccd1 vccd1 _0793_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_23_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1414_ _1415_/A vssd1 vssd1 vccd1 vccd1 _1414_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_3_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1276_ _1384_/A vssd1 vssd1 vccd1 vccd1 _1276_/Y sky130_fd_sc_hd__inv_2
X_1345_ _1384_/A vssd1 vssd1 vccd1 vccd1 _1345_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1046__B2 _1071_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout132 _1324_/A vssd1 vssd1 vccd1 vccd1 _1405_/A sky130_fd_sc_hd__buf_6
Xfanout121 _1416_/A vssd1 vssd1 vccd1 vccd1 _1387_/A sky130_fd_sc_hd__buf_8
XFILLER_0_1_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout110 _0970_/X vssd1 vssd1 vccd1 vccd1 _1103_/B sky130_fd_sc_hd__buf_8
XANTENNA__1037__B2 _1030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1130_ hold154/X hold167/X _1135_/S vssd1 vssd1 vccd1 vccd1 _1130_/X sky130_fd_sc_hd__mux2_1
X_1061_ hold68/X _1061_/A2 _1023_/Y hold165/X vssd1 vssd1 vccd1 vccd1 _1507_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_34_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0914_ _0913_/B _0913_/Y _0914_/S vssd1 vssd1 vccd1 vccd1 _0914_/X sky130_fd_sc_hd__mux2_1
X_0845_ _1606_/Q _0831_/A _0845_/S vssd1 vssd1 vccd1 vccd1 _0845_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1028__B2 _1027_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0776_ _0776_/A _0801_/B vssd1 vssd1 vccd1 vccd1 _0831_/A sky130_fd_sc_hd__and2_2
XFILLER_0_11_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1259_ _1339_/A vssd1 vssd1 vccd1 vccd1 _1259_/Y sky130_fd_sc_hd__inv_2
X_1328_ _1415_/A vssd1 vssd1 vccd1 vccd1 _1328_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_46_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1103__B _1103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0955__A_N _1100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1113_ hold44/X _1478_/Q _1135_/S vssd1 vssd1 vccd1 vccd1 hold45/A sky130_fd_sc_hd__mux2_1
XFILLER_0_45_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1044_ _1021_/A _1031_/Y hold28/X _1071_/S vssd1 vssd1 vccd1 vccd1 _1524_/D sky130_fd_sc_hd__a2bb2o_1
XANTENNA__1013__B _1027_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0759_ _0882_/B _0744_/X _0758_/Y _0757_/X vssd1 vssd1 vccd1 vccd1 _1631_/D sky130_fd_sc_hd__a31o_1
X_0828_ _0828_/A _0836_/A vssd1 vssd1 vccd1 vccd1 _0828_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_fanout111_A _1071_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold207 _1169_/X vssd1 vssd1 vccd1 vccd1 _1428_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold229 _1497_/Q vssd1 vssd1 vccd1 vccd1 _1137_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold218 _1431_/Q vssd1 vssd1 vccd1 vccd1 hold218/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1593_ _1632_/CLK hold5/X _1375_/Y vssd1 vssd1 vccd1 vccd1 _1593_/Q sky130_fd_sc_hd__dfrtp_1
X_1027_ _1027_/A _1027_/B vssd1 vssd1 vccd1 vccd1 _1027_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_56_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1100__C _1100_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0948__A _1100_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold90 hold90/A vssd1 vssd1 vccd1 vccd1 hold90/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1576_ _1580_/CLK _1576_/D _1358_/Y vssd1 vssd1 vccd1 vccd1 _1576_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1430_ _1547_/CLK hold37/X _1212_/Y vssd1 vssd1 vccd1 vccd1 _1430_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput80 _1474_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[18] sky130_fd_sc_hd__buf_12
X_1361_ _1363_/A vssd1 vssd1 vccd1 vccd1 _1361_/Y sky130_fd_sc_hd__inv_2
X_1292_ _1324_/A vssd1 vssd1 vccd1 vccd1 _1292_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput91 _1484_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[28] sky130_fd_sc_hd__buf_12
XFILLER_0_26_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1021__B _1027_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1559_ _1623_/CLK _1559_/D _1341_/Y vssd1 vssd1 vccd1 vccd1 hold44/A sky130_fd_sc_hd__dfrtp_1
X_1628_ _1632_/CLK _1628_/D _1410_/Y vssd1 vssd1 vccd1 vccd1 hold40/A sky130_fd_sc_hd__dfrtp_1
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold390 _1574_/Q vssd1 vssd1 vccd1 vccd1 hold390/X sky130_fd_sc_hd__dlygate4sd3_1
X_0930_ _1568_/Q _1567_/Q _0886_/B vssd1 vssd1 vccd1 vccd1 _0930_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_23_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1055__A2 _1059_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_20_clk_A clkbuf_1_1__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0861_ hold124/X hold141/X _0865_/S vssd1 vssd1 vccd1 vccd1 _0861_/X sky130_fd_sc_hd__mux2_1
X_0792_ _0792_/A vssd1 vssd1 vccd1 vccd1 _1624_/D sky130_fd_sc_hd__inv_2
XFILLER_0_48_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1413_ _1413_/A vssd1 vssd1 vccd1 vccd1 _1413_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_23_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1344_ _1387_/A vssd1 vssd1 vccd1 vccd1 _1344_/Y sky130_fd_sc_hd__inv_2
X_1275_ _1384_/A vssd1 vssd1 vccd1 vccd1 _1275_/Y sky130_fd_sc_hd__inv_2
Xfanout133 _1324_/A vssd1 vssd1 vccd1 vccd1 _1397_/A sky130_fd_sc_hd__buf_8
Xfanout122 _1416_/A vssd1 vssd1 vccd1 vccd1 _1410_/A sky130_fd_sc_hd__buf_4
Xfanout111 _1071_/S vssd1 vssd1 vccd1 vccd1 _1069_/S sky130_fd_sc_hd__buf_4
XFILLER_0_49_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1060_ hold88/X _1069_/S _1021_/Y _1031_/C vssd1 vssd1 vccd1 vccd1 _1060_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_34_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0913_ _0913_/A _0913_/B vssd1 vssd1 vccd1 vccd1 _0913_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0844_ _0782_/X _0793_/Y _0843_/X _0831_/A _0843_/A vssd1 vssd1 vccd1 vccd1 _0844_/X
+ sky130_fd_sc_hd__a32o_1
X_0775_ _0775_/A _1101_/B vssd1 vssd1 vccd1 vccd1 _0801_/B sky130_fd_sc_hd__nand2_1
X_1258_ _1339_/A vssd1 vssd1 vccd1 vccd1 _1258_/Y sky130_fd_sc_hd__inv_2
X_1327_ _1384_/A vssd1 vssd1 vccd1 vccd1 _1327_/Y sky130_fd_sc_hd__inv_2
X_1189_ hold277/X _1187_/X _1188_/X _1185_/A vssd1 vssd1 vccd1 vccd1 _1189_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_19_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1194__A1 _0995_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1112_ hold175/X _1479_/Q _1135_/S vssd1 vssd1 vccd1 vccd1 _1112_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1043_ _1019_/A _1031_/Y hold50/X _1059_/A2 vssd1 vssd1 vccd1 vccd1 _1043_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_43_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0827_ _0833_/A _1613_/Q _0835_/B vssd1 vssd1 vccd1 vccd1 _0829_/S sky130_fd_sc_hd__and3_1
X_0758_ _0764_/D _0758_/B vssd1 vssd1 vccd1 vccd1 _0758_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold208 _1631_/Q vssd1 vssd1 vccd1 vccd1 hold208/X sky130_fd_sc_hd__dlygate4sd3_1
X_1592_ _1634_/CLK hold3/X _1374_/Y vssd1 vssd1 vccd1 vccd1 _1592_/Q sky130_fd_sc_hd__dfrtp_1
Xhold219 _1166_/X vssd1 vssd1 vccd1 vccd1 _1431_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1026_ hold149/X _1071_/S _1103_/B _1025_/Y vssd1 vssd1 vccd1 vccd1 _1026_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_16_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0948__B _1007_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold80 hold80/A vssd1 vssd1 vccd1 vccd1 hold80/X sky130_fd_sc_hd__clkbuf_2
Xhold91 hold91/A vssd1 vssd1 vccd1 vccd1 hold91/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1575_ _1580_/CLK _1575_/D _1357_/Y vssd1 vssd1 vccd1 vccd1 _1575_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1019__B _1027_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1009_ hold90/X _1069_/S _1103_/B _1008_/X vssd1 vssd1 vccd1 vccd1 hold91/A sky130_fd_sc_hd__a22o_1
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1000__B1 _1103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput70 _1636_/A vssd1 vssd1 vccd1 vccd1 wb_cyc_o sky130_fd_sc_hd__buf_12
X_1360_ _1364_/A vssd1 vssd1 vccd1 vccd1 _1360_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_50_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1291_ _1324_/A vssd1 vssd1 vccd1 vccd1 _1291_/Y sky130_fd_sc_hd__inv_2
Xoutput92 _1485_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[29] sky130_fd_sc_hd__buf_12
Xoutput81 _1475_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[19] sky130_fd_sc_hd__buf_12
XFILLER_0_53_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_9_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1489_ _1489_/CLK _1489_/D _1271_/Y vssd1 vssd1 vccd1 vccd1 _1489_/Q sky130_fd_sc_hd__dfrtp_1
X_1627_ _1627_/CLK _1627_/D _1409_/Y vssd1 vssd1 vccd1 vccd1 _1627_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1558_ _1558_/CLK _1558_/D _1340_/Y vssd1 vssd1 vccd1 vccd1 hold66/A sky130_fd_sc_hd__dfrtp_1
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold380 _1591_/Q vssd1 vssd1 vccd1 vccd1 hold380/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_25_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _1605_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_23_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0860_ hold62/X hold104/X _0865_/S vssd1 vssd1 vccd1 vccd1 hold63/A sky130_fd_sc_hd__mux2_1
X_0791_ _0783_/X hold313/X _0851_/S vssd1 vssd1 vccd1 vccd1 _0792_/A sky130_fd_sc_hd__mux2_1
X_1412_ _1413_/A vssd1 vssd1 vccd1 vccd1 _1412_/Y sky130_fd_sc_hd__inv_2
X_1343_ _1387_/A vssd1 vssd1 vccd1 vccd1 _1343_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_3_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1274_ _1385_/A vssd1 vssd1 vccd1 vccd1 _1274_/Y sky130_fd_sc_hd__inv_2
XANTENNA_fanout134_A _1416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_16_clk clkbuf_1_1__f_clk/X vssd1 vssd1 vccd1 vccd1 _1625_/CLK sky130_fd_sc_hd__clkbuf_16
X_0989_ _1100_/A _1007_/B _0989_/C vssd1 vssd1 vccd1 vccd1 _0990_/B sky130_fd_sc_hd__and3b_1
XFILLER_0_14_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout134 _1416_/A vssd1 vssd1 vccd1 vccd1 _1324_/A sky130_fd_sc_hd__buf_4
Xfanout123 _1364_/A vssd1 vssd1 vccd1 vccd1 _1417_/A sky130_fd_sc_hd__buf_8
Xfanout112 _1068_/S vssd1 vssd1 vccd1 vccd1 _1071_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0912_ _0912_/A _0933_/B _0915_/C _0915_/D vssd1 vssd1 vccd1 vccd1 _0913_/B sky130_fd_sc_hd__and4_1
XFILLER_0_34_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0843_ _0843_/A _1608_/Q vssd1 vssd1 vccd1 vccd1 _0843_/X sky130_fd_sc_hd__or2_1
X_0774_ _0776_/A _0774_/B vssd1 vssd1 vccd1 vccd1 _0784_/B sky130_fd_sc_hd__nor2_2
X_1326_ _1405_/A vssd1 vssd1 vccd1 vccd1 _1326_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_5_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _1586_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__1027__B _1027_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1257_ _1339_/A vssd1 vssd1 vccd1 vccd1 _1257_/Y sky130_fd_sc_hd__inv_2
X_1188_ _1136_/B _1136_/D _1188_/C _1188_/D vssd1 vssd1 vccd1 vccd1 _1188_/X sky130_fd_sc_hd__and4bb_1
XFILLER_0_46_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1194__A2 _1007_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1111_ _1192_/C hold306/X _1133_/S vssd1 vssd1 vccd1 vccd1 _1480_/D sky130_fd_sc_hd__mux2_1
X_1042_ _0975_/X _1031_/Y hold42/X _1059_/A2 vssd1 vssd1 vccd1 vccd1 hold87/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0757_ _0753_/A _0726_/A _0753_/D hold208/X vssd1 vssd1 vccd1 vccd1 _0757_/X sky130_fd_sc_hd__o31a_1
X_0826_ _0837_/A _0826_/B _0837_/B vssd1 vssd1 vccd1 vccd1 _0835_/B sky130_fd_sc_hd__and3_1
XFILLER_0_10_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1309_ _1385_/A vssd1 vssd1 vccd1 vccd1 _1309_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_19_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold209 _0871_/X vssd1 vssd1 vccd1 vccd1 _1590_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1591_ _1632_/CLK _1591_/D _1373_/Y vssd1 vssd1 vccd1 vccd1 _1591_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1025_ _1025_/A _1027_/B vssd1 vssd1 vccd1 vccd1 _1025_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_8_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0809_ _0807_/A _0812_/A _0836_/A vssd1 vssd1 vccd1 vccd1 _0810_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_21_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold92 hold92/A vssd1 vssd1 vccd1 vccd1 hold92/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 hold70/A vssd1 vssd1 vccd1 vccd1 hold70/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 hold81/A vssd1 vssd1 vccd1 vccd1 hold81/X sky130_fd_sc_hd__buf_2
XFILLER_0_53_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1574_ _1589_/CLK _1574_/D _1356_/Y vssd1 vssd1 vccd1 vccd1 _1574_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1076__A1 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1008_ hold81/X _1008_/B vssd1 vssd1 vccd1 vccd1 _1008_/X sky130_fd_sc_hd__and2_1
XFILLER_0_50_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput60 _1426_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[2] sky130_fd_sc_hd__buf_12
Xoutput82 _1457_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[1] sky130_fd_sc_hd__buf_12
XFILLER_0_50_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput71 _1456_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[0] sky130_fd_sc_hd__buf_12
Xoutput93 _1458_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[2] sky130_fd_sc_hd__buf_12
XFILLER_0_10_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1290_ _1339_/A vssd1 vssd1 vccd1 vccd1 _1290_/Y sky130_fd_sc_hd__inv_2
XANTENNA__0975__A _1100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1058__B2 _1029_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1626_ _1627_/CLK _1626_/D _1408_/Y vssd1 vssd1 vccd1 vccd1 _1626_/Q sky130_fd_sc_hd__dfrtp_1
X_1488_ _1602_/CLK _1488_/D _1270_/Y vssd1 vssd1 vccd1 vccd1 _1488_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1557_ _1558_/CLK _1557_/D _1339_/Y vssd1 vssd1 vccd1 vccd1 _1557_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1049__B2 _1031_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold381 _1544_/Q vssd1 vssd1 vccd1 vccd1 hold381/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold370 _1587_/Q vssd1 vssd1 vccd1 vccd1 hold370/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0790_ _0767_/Y hold313/X _0789_/X _0783_/X _0789_/A vssd1 vssd1 vccd1 vccd1 _0790_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_2_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1342_ _1404_/A vssd1 vssd1 vccd1 vccd1 _1342_/Y sky130_fd_sc_hd__inv_2
X_1411_ _1413_/A vssd1 vssd1 vccd1 vccd1 _1411_/Y sky130_fd_sc_hd__inv_2
X_1273_ _1402_/A vssd1 vssd1 vccd1 vccd1 _1273_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_3_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout127_A _1416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0988_ hold86/X hold80/X vssd1 vssd1 vccd1 vccd1 _1027_/B sky130_fd_sc_hd__or2_4
X_1609_ _1623_/CLK _1609_/D _1391_/Y vssd1 vssd1 vccd1 vccd1 _1609_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout113 _1059_/A2 vssd1 vssd1 vccd1 vccd1 _1061_/A2 sky130_fd_sc_hd__buf_4
XFILLER_0_1_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout135 input3/X vssd1 vssd1 vccd1 vccd1 _1416_/A sky130_fd_sc_hd__buf_8
Xfanout124 _1364_/A vssd1 vssd1 vccd1 vccd1 _1363_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_52_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_8_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0911_ _0910_/A _0908_/Y _0910_/X vssd1 vssd1 vccd1 vccd1 _0911_/Y sky130_fd_sc_hd__o21bai_1
X_0842_ _0782_/X _0794_/Y _0841_/X _0831_/A _0795_/B vssd1 vssd1 vccd1 vccd1 _0842_/X
+ sky130_fd_sc_hd__a32o_1
X_0773_ _0773_/A _0773_/B _0773_/C _0773_/D vssd1 vssd1 vccd1 vccd1 _0773_/X sky130_fd_sc_hd__or4_1
X_1256_ _1413_/A vssd1 vssd1 vccd1 vccd1 _1256_/Y sky130_fd_sc_hd__inv_2
X_1325_ _1405_/A vssd1 vssd1 vccd1 vccd1 _1325_/Y sky130_fd_sc_hd__inv_2
X_1187_ _1137_/B _1137_/D _1187_/C _1187_/D vssd1 vssd1 vccd1 vccd1 _1187_/X sky130_fd_sc_hd__and4bb_1
XFILLER_0_19_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1110_ _1007_/C hold288/X _1135_/S vssd1 vssd1 vccd1 vccd1 _1481_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_29_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0983__A _1100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1041_ _1015_/A _1031_/Y hold70/X _1059_/A2 vssd1 vssd1 vccd1 vccd1 _1041_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0825_ _0836_/A _0825_/B _0825_/C vssd1 vssd1 vccd1 vccd1 _0825_/X sky130_fd_sc_hd__and3_1
XFILLER_0_28_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0756_ hold24/X _0753_/X _0755_/X vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__a21o_1
XFILLER_0_3_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1239_ _1363_/A vssd1 vssd1 vccd1 vccd1 _1239_/Y sky130_fd_sc_hd__inv_2
X_1308_ _1385_/A vssd1 vssd1 vccd1 vccd1 _1308_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold204_A _1462_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1590_ _1631_/CLK _1590_/D _1372_/Y vssd1 vssd1 vccd1 vccd1 _1590_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1024_ hold64/X _1071_/S _1103_/B _1023_/Y vssd1 vssd1 vccd1 vccd1 hold65/A sky130_fd_sc_hd__a22o_1
XFILLER_0_56_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0808_ _0802_/A _0802_/Y _0808_/S vssd1 vssd1 vccd1 vccd1 _0808_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_12_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0739_ _0739_/A _0896_/A _0919_/A _0923_/S vssd1 vssd1 vccd1 vccd1 _0740_/D sky130_fd_sc_hd__or4b_1
XFILLER_0_39_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1094__A2 input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold93 hold93/A vssd1 vssd1 vccd1 vccd1 hold93/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 hold82/A vssd1 vssd1 vccd1 vccd1 hold82/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 hold60/A vssd1 vssd1 vccd1 vccd1 hold60/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 hold71/A vssd1 vssd1 vccd1 vccd1 hold71/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1085__A2 input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1573_ _1589_/CLK _1573_/D _1355_/Y vssd1 vssd1 vccd1 vccd1 _1573_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1007_ _1564_/Q _1007_/B _1007_/C vssd1 vssd1 vccd1 vccd1 _1007_/X sky130_fd_sc_hd__and3b_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1000__A2 _1071_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput50 _1444_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[20] sky130_fd_sc_hd__buf_12
Xoutput72 _1466_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[10] sky130_fd_sc_hd__buf_12
Xoutput83 _1476_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[20] sky130_fd_sc_hd__buf_12
Xoutput61 _1454_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[30] sky130_fd_sc_hd__buf_12
Xoutput94 _1486_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[30] sky130_fd_sc_hd__buf_12
XFILLER_0_53_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0975__B _1007_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1625_ _1625_/CLK _1625_/D _1407_/Y vssd1 vssd1 vccd1 vccd1 _1625_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1556_ _1556_/CLK hold95/X _1338_/Y vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__dfrtp_1
X_1487_ _1548_/CLK _1487_/D _1269_/Y vssd1 vssd1 vccd1 vccd1 _1487_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_27_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1049__A2 _1069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold360 _1613_/Q vssd1 vssd1 vccd1 vccd1 _0835_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 _1589_/Q vssd1 vssd1 vccd1 vccd1 hold371/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 _1592_/Q vssd1 vssd1 vccd1 vccd1 hold382/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0980__B2 _1069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1410_ _1410_/A vssd1 vssd1 vccd1 vccd1 _1410_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_23_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1341_ _1404_/A vssd1 vssd1 vccd1 vccd1 _1341_/Y sky130_fd_sc_hd__inv_2
X_1272_ _1402_/A vssd1 vssd1 vccd1 vccd1 _1272_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_13_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0987_ _1563_/Q hold80/X vssd1 vssd1 vccd1 vccd1 hold81/A sky130_fd_sc_hd__nor2_1
Xfanout125 _1364_/A vssd1 vssd1 vccd1 vccd1 _1413_/A sky130_fd_sc_hd__buf_8
X_1608_ _1623_/CLK _1608_/D _1390_/Y vssd1 vssd1 vccd1 vccd1 _1608_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout114 _1068_/S vssd1 vssd1 vccd1 vccd1 _1059_/A2 sky130_fd_sc_hd__buf_4
XFILLER_0_1_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1539_ _1605_/CLK hold65/X _1321_/Y vssd1 vssd1 vccd1 vccd1 hold64/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold190 _1584_/Q vssd1 vssd1 vccd1 vccd1 _0764_/A sky130_fd_sc_hd__buf_2
XFILLER_0_34_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0910_ _0910_/A _0933_/B _0910_/C vssd1 vssd1 vccd1 vccd1 _0910_/X sky130_fd_sc_hd__and3_1
X_0841_ _1609_/Q _1608_/Q _0795_/B vssd1 vssd1 vccd1 vccd1 _0841_/X sky130_fd_sc_hd__a21o_1
X_0772_ _1617_/Q _1616_/Q _1615_/Q _0833_/A vssd1 vssd1 vccd1 vccd1 _0773_/D sky130_fd_sc_hd__or4b_1
XFILLER_0_11_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1255_ _1363_/A vssd1 vssd1 vccd1 vccd1 _1255_/Y sky130_fd_sc_hd__inv_2
X_1324_ _1324_/A vssd1 vssd1 vccd1 vccd1 _1324_/Y sky130_fd_sc_hd__inv_2
X_1186_ _1183_/Y _1185_/X _1179_/A _1179_/B vssd1 vssd1 vccd1 vccd1 _1420_/D sky130_fd_sc_hd__a211o_1
XFILLER_0_46_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1340__A _1416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0871__A0 hold84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1040_ _1013_/A _1031_/Y hold239/X _1061_/A2 vssd1 vssd1 vccd1 vccd1 _1528_/D sky130_fd_sc_hd__a2bb2o_1
XANTENNA__0983__B _1007_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0824_ _0837_/A _1606_/Q _0837_/B _0804_/C _0803_/D vssd1 vssd1 vccd1 vccd1 _0824_/X
+ sky130_fd_sc_hd__a41o_1
X_0755_ _0753_/D _0755_/B vssd1 vssd1 vccd1 vccd1 _0755_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1169_ hold195/X hold206/X _1171_/S vssd1 vssd1 vccd1 vccd1 _1169_/X sky130_fd_sc_hd__mux2_1
X_1307_ _1324_/A vssd1 vssd1 vccd1 vccd1 _1307_/Y sky130_fd_sc_hd__inv_2
X_1238_ _1404_/A vssd1 vssd1 vccd1 vccd1 _1238_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_7_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1097__A0 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1023_ _1023_/A _1027_/B vssd1 vssd1 vccd1 vccd1 _1023_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__1088__A0 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0738_ _0886_/A _0886_/C _1567_/Q _0886_/B vssd1 vssd1 vccd1 vccd1 _0740_/C sky130_fd_sc_hd__or4bb_1
X_0807_ _0807_/A _0812_/A vssd1 vssd1 vccd1 vccd1 _0808_/S sky130_fd_sc_hd__nand2_1
XFILLER_0_31_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1012__B1 _1103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1079__A0 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1003__B1 _1103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold50 hold50/A vssd1 vssd1 vccd1 vccd1 hold50/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 hold72/A vssd1 vssd1 vccd1 vccd1 hold72/X sky130_fd_sc_hd__buf_1
Xhold83 hold83/A vssd1 vssd1 vccd1 vccd1 hold83/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 hold61/A vssd1 vssd1 vccd1 vccd1 hold61/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 hold94/A vssd1 vssd1 vccd1 vccd1 hold94/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1572_ _1589_/CLK _1572_/D _1354_/Y vssd1 vssd1 vccd1 vccd1 _1572_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1006_ hold156/X _1059_/A2 _1103_/B _1005_/X vssd1 vssd1 vccd1 vccd1 _1006_/X sky130_fd_sc_hd__a22o_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput73 _1467_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[11] sky130_fd_sc_hd__buf_12
Xoutput40 _1435_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[11] sky130_fd_sc_hd__buf_12
Xoutput95 _1487_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[31] sky130_fd_sc_hd__buf_12
Xoutput84 _1477_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[21] sky130_fd_sc_hd__buf_12
Xoutput51 _1445_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[21] sky130_fd_sc_hd__buf_12
Xoutput62 _1455_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[31] sky130_fd_sc_hd__buf_12
XFILLER_0_26_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1555_ _1589_/CLK _1555_/D _1337_/Y vssd1 vssd1 vccd1 vccd1 _1555_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1624_ _1624_/CLK _1624_/D _1406_/Y vssd1 vssd1 vccd1 vccd1 _1624_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1486_ _1605_/CLK _1486_/D _1268_/Y vssd1 vssd1 vccd1 vccd1 _1486_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_19_clk clkbuf_1_1__f_clk/X vssd1 vssd1 vccd1 vccd1 _1547_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold383 _1534_/Q vssd1 vssd1 vccd1 vccd1 hold383/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 _1571_/Q vssd1 vssd1 vccd1 vccd1 _0737_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold350 _1608_/Q vssd1 vssd1 vccd1 vccd1 _0845_/S sky130_fd_sc_hd__dlygate4sd3_1
Xhold372 _1589_/Q vssd1 vssd1 vccd1 vccd1 hold372/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1340_ _1416_/A vssd1 vssd1 vccd1 vccd1 _1340_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_48_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1271_ _1402_/A vssd1 vssd1 vccd1 vccd1 _1271_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_13_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_8_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _1580_/CLK sky130_fd_sc_hd__clkbuf_16
X_0986_ _0971_/Y hold118/X hold10/X _1059_/A2 vssd1 vssd1 vccd1 vccd1 _0986_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_13_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout126 _1416_/A vssd1 vssd1 vccd1 vccd1 _1364_/A sky130_fd_sc_hd__clkbuf_8
X_1469_ _1580_/CLK hold53/X _1251_/Y vssd1 vssd1 vccd1 vccd1 _1469_/Q sky130_fd_sc_hd__dfrtp_2
X_1538_ _1583_/CLK _1538_/D _1320_/Y vssd1 vssd1 vccd1 vccd1 _1538_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1607_ _1625_/CLK _1607_/D _1389_/Y vssd1 vssd1 vccd1 vccd1 _1607_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_1_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout115 _0981_/A vssd1 vssd1 vccd1 vccd1 _1100_/A sky130_fd_sc_hd__buf_4
XFILLER_0_54_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold180 _1545_/Q vssd1 vssd1 vccd1 vccd1 hold180/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold191 _0764_/X vssd1 vssd1 vccd1 vccd1 _0765_/S sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0840_ _1606_/Q _0796_/Y _0839_/X _0831_/A _0795_/A vssd1 vssd1 vccd1 vccd1 _0840_/X
+ sky130_fd_sc_hd__a32o_1
X_0771_ _1613_/Q _1612_/Q _0795_/A _1609_/Q vssd1 vssd1 vccd1 vccd1 _0773_/C sky130_fd_sc_hd__or4_1
X_1323_ _1324_/A vssd1 vssd1 vccd1 vccd1 _1323_/Y sky130_fd_sc_hd__inv_2
X_1254_ _1384_/A vssd1 vssd1 vccd1 vccd1 _1254_/Y sky130_fd_sc_hd__inv_2
X_1185_ _1185_/A _1185_/B _1185_/C vssd1 vssd1 vccd1 vccd1 _1185_/X sky130_fd_sc_hd__or3_1
XFILLER_0_46_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0969_ _1191_/A _0981_/A _1007_/B vssd1 vssd1 vccd1 vccd1 _1013_/A sky130_fd_sc_hd__or3_1
XFILLER_0_6_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0754_ _0754_/A _1583_/Q hold30/A _0764_/C vssd1 vssd1 vccd1 vccd1 _0755_/B sky130_fd_sc_hd__and4_1
X_0823_ _0825_/B hold338/X _0816_/X vssd1 vssd1 vccd1 vccd1 _0823_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1306_ _1417_/A vssd1 vssd1 vccd1 vccd1 _1306_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_19_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1168_ hold158/X hold184/X _1168_/S vssd1 vssd1 vccd1 vccd1 _1168_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_35_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1099_ _1098_/X hold8/X _1099_/S vssd1 vssd1 vccd1 vccd1 _1489_/D sky130_fd_sc_hd__mux2_1
X_1237_ _1339_/A vssd1 vssd1 vccd1 vccd1 _1237_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_42_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1022_ hold230/X _1069_/S _1103_/B _1021_/Y vssd1 vssd1 vccd1 vccd1 _1540_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1088__A1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1110__S _1135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0737_ _0914_/S _0912_/A _0889_/C _0737_/D vssd1 vssd1 vccd1 vccd1 _0740_/B sky130_fd_sc_hd__or4_1
X_0806_ _0806_/A _0813_/A _0826_/B _0813_/B vssd1 vssd1 vccd1 vccd1 _0812_/A sky130_fd_sc_hd__and4_1
XFILLER_0_24_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A vssd1 vssd1 vccd1 vccd1 hold51/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 hold84/A vssd1 vssd1 vccd1 vccd1 hold84/X sky130_fd_sc_hd__clkbuf_2
Xhold73 hold73/A vssd1 vssd1 vccd1 vccd1 hold73/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 hold95/A vssd1 vssd1 vccd1 vccd1 hold95/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 hold62/A vssd1 vssd1 vccd1 vccd1 hold62/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1571_ _1589_/CLK _1571_/D _1353_/Y vssd1 vssd1 vccd1 vccd1 _1571_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0989__B _1007_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_6_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1105__S _1133_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1005_ hold81/X _1005_/B vssd1 vssd1 vccd1 vccd1 _1005_/X sky130_fd_sc_hd__and2_1
XFILLER_0_12_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput52 _1446_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[22] sky130_fd_sc_hd__buf_12
Xoutput41 _1436_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[12] sky130_fd_sc_hd__buf_12
Xoutput85 _1478_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[22] sky130_fd_sc_hd__buf_12
Xoutput96 _1459_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[3] sky130_fd_sc_hd__buf_12
Xoutput74 _1468_/Q vssd1 vssd1 vccd1 vccd1 wb_dat_o[12] sky130_fd_sc_hd__buf_12
Xoutput63 _1427_/Q vssd1 vssd1 vccd1 vccd1 wb_adr_o[3] sky130_fd_sc_hd__buf_12
XFILLER_0_26_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1554_ _1586_/CLK _1554_/D _1336_/Y vssd1 vssd1 vccd1 vccd1 _1554_/Q sky130_fd_sc_hd__dfrtp_1
X_1623_ _1623_/CLK _1623_/D _1405_/Y vssd1 vssd1 vccd1 vccd1 _1623_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1485_ _1556_/CLK _1485_/D _1267_/Y vssd1 vssd1 vccd1 vccd1 _1485_/Q sky130_fd_sc_hd__dfrtp_1
.ends

