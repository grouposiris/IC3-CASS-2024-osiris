magic
tech sky130A
magscale 1 2
timestamp 1730916576
<< nwell >>
rect 1066 2159 148894 127313
<< obsli1 >>
rect 1104 2159 148856 127313
<< obsm1 >>
rect 842 484 148856 129600
<< metal2 >>
rect 18694 129200 18750 130000
rect 19338 129200 19394 130000
rect 19982 129200 20038 130000
rect 20626 129200 20682 130000
rect 74722 129200 74778 130000
rect 75366 129200 75422 130000
rect 76010 129200 76066 130000
rect 76654 129200 76710 130000
rect 77298 129200 77354 130000
rect 77942 129200 77998 130000
rect 78586 129200 78642 130000
rect 79230 129200 79286 130000
rect 79874 129200 79930 130000
rect 80518 129200 80574 130000
rect 81162 129200 81218 130000
rect 81806 129200 81862 130000
rect 82450 129200 82506 130000
rect 83094 129200 83150 130000
rect 85026 129200 85082 130000
rect 85670 129200 85726 130000
rect 86314 129200 86370 130000
rect 86958 129200 87014 130000
rect 87602 129200 87658 130000
rect 137190 129200 137246 130000
rect 137834 129200 137890 130000
rect 138478 129200 138534 130000
rect 139122 129200 139178 130000
rect 141698 129200 141754 130000
rect 142342 129200 142398 130000
rect 142986 129200 143042 130000
rect 143630 129200 143686 130000
rect 4526 0 4582 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 73434 0 73490 800
rect 74722 0 74778 800
rect 75366 0 75422 800
rect 76010 0 76066 800
rect 76654 0 76710 800
rect 79874 0 79930 800
rect 80518 0 80574 800
rect 81162 0 81218 800
rect 81806 0 81862 800
rect 82450 0 82506 800
rect 83094 0 83150 800
rect 85026 0 85082 800
rect 85670 0 85726 800
rect 86314 0 86370 800
rect 86958 0 87014 800
rect 87602 0 87658 800
rect 88246 0 88302 800
<< obsm2 >>
rect 846 129144 18638 129713
rect 18806 129144 19282 129713
rect 19450 129144 19926 129713
rect 20094 129144 20570 129713
rect 20738 129144 74666 129713
rect 74834 129144 75310 129713
rect 75478 129144 75954 129713
rect 76122 129144 76598 129713
rect 76766 129144 77242 129713
rect 77410 129144 77886 129713
rect 78054 129144 78530 129713
rect 78698 129144 79174 129713
rect 79342 129144 79818 129713
rect 79986 129144 80462 129713
rect 80630 129144 81106 129713
rect 81274 129144 81750 129713
rect 81918 129144 82394 129713
rect 82562 129144 83038 129713
rect 83206 129144 84970 129713
rect 85138 129144 85614 129713
rect 85782 129144 86258 129713
rect 86426 129144 86902 129713
rect 87070 129144 87546 129713
rect 87714 129144 137134 129713
rect 137302 129144 137778 129713
rect 137946 129144 138422 129713
rect 138590 129144 139066 129713
rect 139234 129144 141642 129713
rect 141810 129144 142286 129713
rect 142454 129144 142930 129713
rect 143098 129144 143574 129713
rect 143742 129144 148836 129713
rect 846 856 148836 129144
rect 846 439 4470 856
rect 4638 439 6402 856
rect 6570 439 7046 856
rect 7214 439 7690 856
rect 7858 439 8334 856
rect 8502 439 10910 856
rect 11078 439 11554 856
rect 11722 439 12198 856
rect 12366 439 12842 856
rect 13010 439 73378 856
rect 73546 439 74666 856
rect 74834 439 75310 856
rect 75478 439 75954 856
rect 76122 439 76598 856
rect 76766 439 79818 856
rect 79986 439 80462 856
rect 80630 439 81106 856
rect 81274 439 81750 856
rect 81918 439 82394 856
rect 82562 439 83038 856
rect 83206 439 84970 856
rect 85138 439 85614 856
rect 85782 439 86258 856
rect 86426 439 86902 856
rect 87070 439 87546 856
rect 87714 439 88190 856
rect 88358 439 148836 856
<< metal3 >>
rect 149200 82968 150000 83088
rect 149200 82288 150000 82408
rect 149200 81608 150000 81728
rect 149200 80928 150000 81048
rect 0 79568 800 79688
rect 149200 70048 150000 70168
rect 149200 67328 150000 67448
rect 149200 66648 150000 66768
rect 149200 65968 150000 66088
rect 0 65288 800 65408
rect 149200 65288 150000 65408
rect 0 64608 800 64728
rect 149200 64608 150000 64728
rect 149200 61208 150000 61328
rect 149200 59168 150000 59288
rect 149200 51008 150000 51128
rect 0 50328 800 50448
rect 149200 50328 150000 50448
rect 0 49648 800 49768
rect 0 48968 800 49088
rect 149200 35368 150000 35488
rect 149200 30608 150000 30728
rect 149200 24488 150000 24608
<< obsm3 >>
rect 798 83168 149200 129709
rect 798 82888 149120 83168
rect 798 82488 149200 82888
rect 798 82208 149120 82488
rect 798 81808 149200 82208
rect 798 81528 149120 81808
rect 798 81128 149200 81528
rect 798 80848 149120 81128
rect 798 79768 149200 80848
rect 880 79488 149200 79768
rect 798 70248 149200 79488
rect 798 69968 149120 70248
rect 798 67528 149200 69968
rect 798 67248 149120 67528
rect 798 66848 149200 67248
rect 798 66568 149120 66848
rect 798 66168 149200 66568
rect 798 65888 149120 66168
rect 798 65488 149200 65888
rect 880 65208 149120 65488
rect 798 64808 149200 65208
rect 880 64528 149120 64808
rect 798 61408 149200 64528
rect 798 61128 149120 61408
rect 798 59368 149200 61128
rect 798 59088 149120 59368
rect 798 51208 149200 59088
rect 798 50928 149120 51208
rect 798 50528 149200 50928
rect 880 50248 149120 50528
rect 798 49848 149200 50248
rect 880 49568 149200 49848
rect 798 49168 149200 49568
rect 880 48888 149200 49168
rect 798 35568 149200 48888
rect 798 35288 149120 35568
rect 798 30808 149200 35288
rect 798 30528 149120 30808
rect 798 24688 149200 30528
rect 798 24408 149120 24688
rect 798 443 149200 24408
<< metal4 >>
rect 4208 2128 4528 127344
rect 4868 2128 5188 127344
rect 40208 2128 40528 127344
rect 40868 2128 41188 127344
rect 76208 2128 76528 127344
rect 76868 2128 77188 127344
rect 112208 2128 112528 127344
rect 112868 2128 113188 127344
rect 148208 2128 148528 127344
<< obsm4 >>
rect 5395 127424 146957 129709
rect 5395 2048 40128 127424
rect 40608 2048 40788 127424
rect 41268 2048 76128 127424
rect 76608 2048 76788 127424
rect 77268 2048 112128 127424
rect 112608 2048 112788 127424
rect 113268 2048 146957 127424
rect 5395 443 146957 2048
<< labels >>
rlabel metal2 s 4526 0 4582 800 6 clk
port 1 nsew signal input
rlabel metal3 s 149200 70048 150000 70168 6 funct3[0]
port 2 nsew signal input
rlabel metal3 s 149200 30608 150000 30728 6 funct3[1]
port 3 nsew signal input
rlabel metal3 s 149200 65288 150000 65408 6 funct3[2]
port 4 nsew signal input
rlabel metal3 s 149200 24488 150000 24608 6 rst
port 5 nsew signal input
rlabel metal4 s 4208 2128 4528 127344 6 vccd1
port 6 nsew power bidirectional
rlabel metal4 s 40208 2128 40528 127344 6 vccd1
port 6 nsew power bidirectional
rlabel metal4 s 76208 2128 76528 127344 6 vccd1
port 6 nsew power bidirectional
rlabel metal4 s 112208 2128 112528 127344 6 vccd1
port 6 nsew power bidirectional
rlabel metal4 s 148208 2128 148528 127344 6 vccd1
port 6 nsew power bidirectional
rlabel metal4 s 4868 2128 5188 127344 6 vssd1
port 7 nsew ground bidirectional
rlabel metal4 s 40868 2128 41188 127344 6 vssd1
port 7 nsew ground bidirectional
rlabel metal4 s 76868 2128 77188 127344 6 vssd1
port 7 nsew ground bidirectional
rlabel metal4 s 112868 2128 113188 127344 6 vssd1
port 7 nsew ground bidirectional
rlabel metal2 s 82450 0 82506 800 6 wb_ack_o
port 8 nsew signal output
rlabel metal2 s 18694 129200 18750 130000 6 wb_adr_i[0]
port 9 nsew signal input
rlabel metal2 s 20626 129200 20682 130000 6 wb_adr_i[1]
port 10 nsew signal input
rlabel metal2 s 19338 129200 19394 130000 6 wb_adr_i[2]
port 11 nsew signal input
rlabel metal2 s 19982 129200 20038 130000 6 wb_adr_i[3]
port 12 nsew signal input
rlabel metal2 s 76654 129200 76710 130000 6 wb_adr_i[4]
port 13 nsew signal input
rlabel metal2 s 77298 129200 77354 130000 6 wb_adr_i[5]
port 14 nsew signal input
rlabel metal2 s 77942 129200 77998 130000 6 wb_adr_i[6]
port 15 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 wb_cyc_i
port 16 nsew signal input
rlabel metal2 s 139122 129200 139178 130000 6 wb_dat_i[0]
port 17 nsew signal input
rlabel metal3 s 149200 50328 150000 50448 6 wb_dat_i[10]
port 18 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wb_dat_i[11]
port 19 nsew signal input
rlabel metal2 s 142986 129200 143042 130000 6 wb_dat_i[12]
port 20 nsew signal input
rlabel metal3 s 0 50328 800 50448 6 wb_dat_i[13]
port 21 nsew signal input
rlabel metal3 s 149200 80928 150000 81048 6 wb_dat_i[14]
port 22 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 wb_dat_i[15]
port 23 nsew signal input
rlabel metal2 s 138478 129200 138534 130000 6 wb_dat_i[16]
port 24 nsew signal input
rlabel metal3 s 0 79568 800 79688 6 wb_dat_i[17]
port 25 nsew signal input
rlabel metal3 s 0 65288 800 65408 6 wb_dat_i[18]
port 26 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wb_dat_i[19]
port 27 nsew signal input
rlabel metal3 s 149200 65968 150000 66088 6 wb_dat_i[1]
port 28 nsew signal input
rlabel metal2 s 142342 129200 142398 130000 6 wb_dat_i[20]
port 29 nsew signal input
rlabel metal3 s 0 49648 800 49768 6 wb_dat_i[21]
port 30 nsew signal input
rlabel metal3 s 149200 81608 150000 81728 6 wb_dat_i[22]
port 31 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 wb_dat_i[23]
port 32 nsew signal input
rlabel metal2 s 137834 129200 137890 130000 6 wb_dat_i[24]
port 33 nsew signal input
rlabel metal3 s 149200 66648 150000 66768 6 wb_dat_i[25]
port 34 nsew signal input
rlabel metal3 s 0 64608 800 64728 6 wb_dat_i[26]
port 35 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wb_dat_i[27]
port 36 nsew signal input
rlabel metal2 s 141698 129200 141754 130000 6 wb_dat_i[28]
port 37 nsew signal input
rlabel metal3 s 0 48968 800 49088 6 wb_dat_i[29]
port 38 nsew signal input
rlabel metal3 s 149200 51008 150000 51128 6 wb_dat_i[2]
port 39 nsew signal input
rlabel metal3 s 149200 82288 150000 82408 6 wb_dat_i[30]
port 40 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 wb_dat_i[31]
port 41 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 wb_dat_i[3]
port 42 nsew signal input
rlabel metal2 s 143630 129200 143686 130000 6 wb_dat_i[4]
port 43 nsew signal input
rlabel metal3 s 149200 35368 150000 35488 6 wb_dat_i[5]
port 44 nsew signal input
rlabel metal3 s 149200 82968 150000 83088 6 wb_dat_i[6]
port 45 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 wb_dat_i[7]
port 46 nsew signal input
rlabel metal2 s 137190 129200 137246 130000 6 wb_dat_i[8]
port 47 nsew signal input
rlabel metal3 s 149200 67328 150000 67448 6 wb_dat_i[9]
port 48 nsew signal input
rlabel metal2 s 85026 129200 85082 130000 6 wb_dat_o[0]
port 49 nsew signal output
rlabel metal3 s 149200 61208 150000 61328 6 wb_dat_o[10]
port 50 nsew signal output
rlabel metal2 s 79874 0 79930 800 6 wb_dat_o[11]
port 51 nsew signal output
rlabel metal2 s 79874 129200 79930 130000 6 wb_dat_o[12]
port 52 nsew signal output
rlabel metal2 s 83094 0 83150 800 6 wb_dat_o[13]
port 53 nsew signal output
rlabel metal2 s 81806 129200 81862 130000 6 wb_dat_o[14]
port 54 nsew signal output
rlabel metal2 s 86314 0 86370 800 6 wb_dat_o[15]
port 55 nsew signal output
rlabel metal2 s 87602 129200 87658 130000 6 wb_dat_o[16]
port 56 nsew signal output
rlabel metal2 s 83094 129200 83150 130000 6 wb_dat_o[17]
port 57 nsew signal output
rlabel metal3 s 149200 64608 150000 64728 6 wb_dat_o[18]
port 58 nsew signal output
rlabel metal2 s 75366 0 75422 800 6 wb_dat_o[19]
port 59 nsew signal output
rlabel metal2 s 78586 129200 78642 130000 6 wb_dat_o[1]
port 60 nsew signal output
rlabel metal2 s 76010 129200 76066 130000 6 wb_dat_o[20]
port 61 nsew signal output
rlabel metal2 s 87602 0 87658 800 6 wb_dat_o[21]
port 62 nsew signal output
rlabel metal2 s 85670 129200 85726 130000 6 wb_dat_o[22]
port 63 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 wb_dat_o[23]
port 64 nsew signal output
rlabel metal2 s 86314 129200 86370 130000 6 wb_dat_o[24]
port 65 nsew signal output
rlabel metal2 s 79230 129200 79286 130000 6 wb_dat_o[25]
port 66 nsew signal output
rlabel metal2 s 74722 0 74778 800 6 wb_dat_o[26]
port 67 nsew signal output
rlabel metal2 s 76010 0 76066 800 6 wb_dat_o[27]
port 68 nsew signal output
rlabel metal2 s 75366 129200 75422 130000 6 wb_dat_o[28]
port 69 nsew signal output
rlabel metal2 s 86958 0 87014 800 6 wb_dat_o[29]
port 70 nsew signal output
rlabel metal3 s 149200 59168 150000 59288 6 wb_dat_o[2]
port 71 nsew signal output
rlabel metal2 s 86958 129200 87014 130000 6 wb_dat_o[30]
port 72 nsew signal output
rlabel metal2 s 88246 0 88302 800 6 wb_dat_o[31]
port 73 nsew signal output
rlabel metal2 s 73434 0 73490 800 6 wb_dat_o[3]
port 74 nsew signal output
rlabel metal2 s 74722 129200 74778 130000 6 wb_dat_o[4]
port 75 nsew signal output
rlabel metal2 s 76654 0 76710 800 6 wb_dat_o[5]
port 76 nsew signal output
rlabel metal2 s 80518 129200 80574 130000 6 wb_dat_o[6]
port 77 nsew signal output
rlabel metal2 s 85026 0 85082 800 6 wb_dat_o[7]
port 78 nsew signal output
rlabel metal2 s 82450 129200 82506 130000 6 wb_dat_o[8]
port 79 nsew signal output
rlabel metal2 s 81162 129200 81218 130000 6 wb_dat_o[9]
port 80 nsew signal output
rlabel metal2 s 80518 0 80574 800 6 wb_stb_i
port 81 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 wb_we_i
port 82 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 150000 130000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 80706890
string GDS_FILE /openlane/designs/mem_byte/runs/small/results/signoff/mem_byte.magic.gds
string GDS_START 729100
<< end >>

